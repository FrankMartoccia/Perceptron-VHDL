library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LUT_4096 is
	port (
		address : in  std_logic_vector(11 downto 0);
		sigmoid_out : out std_logic_vector(15 downto 0) 
	);
end LUT_4096;

architecture beh of LUT_4096 is
	type LUT_t is array (natural range 0 to 4095) of integer;
	constant LUT: LUT_t := (
		0 => 16384,
		1 => 16416,
		2 => 16448,
		3 => 16480,
		4 => 16512,
		5 => 16544,
		6 => 16576,
		7 => 16608,
		8 => 16640,
		9 => 16672,
		10 => 16704,
		11 => 16736,
		12 => 16768,
		13 => 16799,
		14 => 16831,
		15 => 16863,
		16 => 16895,
		17 => 16927,
		18 => 16959,
		19 => 16991,
		20 => 17023,
		21 => 17055,
		22 => 17087,
		23 => 17119,
		24 => 17151,
		25 => 17183,
		26 => 17215,
		27 => 17247,
		28 => 17279,
		29 => 17311,
		30 => 17343,
		31 => 17375,
		32 => 17406,
		33 => 17438,
		34 => 17470,
		35 => 17502,
		36 => 17534,
		37 => 17566,
		38 => 17598,
		39 => 17629,
		40 => 17661,
		41 => 17693,
		42 => 17725,
		43 => 17757,
		44 => 17788,
		45 => 17820,
		46 => 17852,
		47 => 17884,
		48 => 17915,
		49 => 17947,
		50 => 17979,
		51 => 18010,
		52 => 18042,
		53 => 18074,
		54 => 18105,
		55 => 18137,
		56 => 18169,
		57 => 18200,
		58 => 18232,
		59 => 18264,
		60 => 18295,
		61 => 18327,
		62 => 18358,
		63 => 18390,
		64 => 18421,
		65 => 18453,
		66 => 18484,
		67 => 18516,
		68 => 18547,
		69 => 18579,
		70 => 18610,
		71 => 18642,
		72 => 18673,
		73 => 18704,
		74 => 18736,
		75 => 18767,
		76 => 18798,
		77 => 18830,
		78 => 18861,
		79 => 18892,
		80 => 18923,
		81 => 18955,
		82 => 18986,
		83 => 19017,
		84 => 19048,
		85 => 19079,
		86 => 19110,
		87 => 19142,
		88 => 19173,
		89 => 19204,
		90 => 19235,
		91 => 19266,
		92 => 19297,
		93 => 19328,
		94 => 19359,
		95 => 19390,
		96 => 19421,
		97 => 19452,
		98 => 19482,
		99 => 19513,
		100 => 19544,
		101 => 19575,
		102 => 19606,
		103 => 19636,
		104 => 19667,
		105 => 19698,
		106 => 19729,
		107 => 19759,
		108 => 19790,
		109 => 19820,
		110 => 19851,
		111 => 19882,
		112 => 19912,
		113 => 19943,
		114 => 19973,
		115 => 20004,
		116 => 20034,
		117 => 20064,
		118 => 20095,
		119 => 20125,
		120 => 20155,
		121 => 20186,
		122 => 20216,
		123 => 20246,
		124 => 20276,
		125 => 20307,
		126 => 20337,
		127 => 20367,
		128 => 20397,
		129 => 20427,
		130 => 20457,
		131 => 20487,
		132 => 20517,
		133 => 20547,
		134 => 20577,
		135 => 20607,
		136 => 20637,
		137 => 20667,
		138 => 20696,
		139 => 20726,
		140 => 20756,
		141 => 20786,
		142 => 20815,
		143 => 20845,
		144 => 20875,
		145 => 20904,
		146 => 20934,
		147 => 20963,
		148 => 20993,
		149 => 21022,
		150 => 21052,
		151 => 21081,
		152 => 21110,
		153 => 21140,
		154 => 21169,
		155 => 21198,
		156 => 21228,
		157 => 21257,
		158 => 21286,
		159 => 21315,
		160 => 21344,
		161 => 21373,
		162 => 21402,
		163 => 21431,
		164 => 21460,
		165 => 21489,
		166 => 21518,
		167 => 21547,
		168 => 21576,
		169 => 21604,
		170 => 21633,
		171 => 21662,
		172 => 21690,
		173 => 21719,
		174 => 21748,
		175 => 21776,
		176 => 21805,
		177 => 21833,
		178 => 21862,
		179 => 21890,
		180 => 21918,
		181 => 21947,
		182 => 21975,
		183 => 22003,
		184 => 22032,
		185 => 22060,
		186 => 22088,
		187 => 22116,
		188 => 22144,
		189 => 22172,
		190 => 22200,
		191 => 22228,
		192 => 22256,
		193 => 22284,
		194 => 22312,
		195 => 22339,
		196 => 22367,
		197 => 22395,
		198 => 22423,
		199 => 22450,
		200 => 22478,
		201 => 22505,
		202 => 22533,
		203 => 22560,
		204 => 22588,
		205 => 22615,
		206 => 22643,
		207 => 22670,
		208 => 22697,
		209 => 22724,
		210 => 22752,
		211 => 22779,
		212 => 22806,
		213 => 22833,
		214 => 22860,
		215 => 22887,
		216 => 22914,
		217 => 22941,
		218 => 22968,
		219 => 22994,
		220 => 23021,
		221 => 23048,
		222 => 23075,
		223 => 23101,
		224 => 23128,
		225 => 23154,
		226 => 23181,
		227 => 23207,
		228 => 23234,
		229 => 23260,
		230 => 23287,
		231 => 23313,
		232 => 23339,
		233 => 23365,
		234 => 23392,
		235 => 23418,
		236 => 23444,
		237 => 23470,
		238 => 23496,
		239 => 23522,
		240 => 23548,
		241 => 23574,
		242 => 23599,
		243 => 23625,
		244 => 23651,
		245 => 23677,
		246 => 23702,
		247 => 23728,
		248 => 23753,
		249 => 23779,
		250 => 23804,
		251 => 23830,
		252 => 23855,
		253 => 23880,
		254 => 23906,
		255 => 23931,
		256 => 23956,
		257 => 23981,
		258 => 24006,
		259 => 24031,
		260 => 24056,
		261 => 24081,
		262 => 24106,
		263 => 24131,
		264 => 24156,
		265 => 24181,
		266 => 24206,
		267 => 24230,
		268 => 24255,
		269 => 24279,
		270 => 24304,
		271 => 24329,
		272 => 24353,
		273 => 24377,
		274 => 24402,
		275 => 24426,
		276 => 24450,
		277 => 24475,
		278 => 24499,
		279 => 24523,
		280 => 24547,
		281 => 24571,
		282 => 24595,
		283 => 24619,
		284 => 24643,
		285 => 24667,
		286 => 24691,
		287 => 24714,
		288 => 24738,
		289 => 24762,
		290 => 24785,
		291 => 24809,
		292 => 24832,
		293 => 24856,
		294 => 24879,
		295 => 24903,
		296 => 24926,
		297 => 24949,
		298 => 24972,
		299 => 24996,
		300 => 25019,
		301 => 25042,
		302 => 25065,
		303 => 25088,
		304 => 25111,
		305 => 25134,
		306 => 25157,
		307 => 25179,
		308 => 25202,
		309 => 25225,
		310 => 25248,
		311 => 25270,
		312 => 25293,
		313 => 25315,
		314 => 25338,
		315 => 25360,
		316 => 25382,
		317 => 25405,
		318 => 25427,
		319 => 25449,
		320 => 25472,
		321 => 25494,
		322 => 25516,
		323 => 25538,
		324 => 25560,
		325 => 25582,
		326 => 25604,
		327 => 25625,
		328 => 25647,
		329 => 25669,
		330 => 25691,
		331 => 25712,
		332 => 25734,
		333 => 25756,
		334 => 25777,
		335 => 25798,
		336 => 25820,
		337 => 25841,
		338 => 25863,
		339 => 25884,
		340 => 25905,
		341 => 25926,
		342 => 25947,
		343 => 25968,
		344 => 25989,
		345 => 26010,
		346 => 26031,
		347 => 26052,
		348 => 26073,
		349 => 26094,
		350 => 26115,
		351 => 26135,
		352 => 26156,
		353 => 26177,
		354 => 26197,
		355 => 26218,
		356 => 26238,
		357 => 26258,
		358 => 26279,
		359 => 26299,
		360 => 26319,
		361 => 26340,
		362 => 26360,
		363 => 26380,
		364 => 26400,
		365 => 26420,
		366 => 26440,
		367 => 26460,
		368 => 26480,
		369 => 26500,
		370 => 26519,
		371 => 26539,
		372 => 26559,
		373 => 26578,
		374 => 26598,
		375 => 26618,
		376 => 26637,
		377 => 26656,
		378 => 26676,
		379 => 26695,
		380 => 26715,
		381 => 26734,
		382 => 26753,
		383 => 26772,
		384 => 26791,
		385 => 26810,
		386 => 26829,
		387 => 26848,
		388 => 26867,
		389 => 26886,
		390 => 26905,
		391 => 26924,
		392 => 26942,
		393 => 26961,
		394 => 26980,
		395 => 26998,
		396 => 27017,
		397 => 27035,
		398 => 27054,
		399 => 27072,
		400 => 27091,
		401 => 27109,
		402 => 27127,
		403 => 27145,
		404 => 27164,
		405 => 27182,
		406 => 27200,
		407 => 27218,
		408 => 27236,
		409 => 27254,
		410 => 27272,
		411 => 27290,
		412 => 27307,
		413 => 27325,
		414 => 27343,
		415 => 27360,
		416 => 27378,
		417 => 27396,
		418 => 27413,
		419 => 27431,
		420 => 27448,
		421 => 27465,
		422 => 27483,
		423 => 27500,
		424 => 27517,
		425 => 27535,
		426 => 27552,
		427 => 27569,
		428 => 27586,
		429 => 27603,
		430 => 27620,
		431 => 27637,
		432 => 27654,
		433 => 27671,
		434 => 27687,
		435 => 27704,
		436 => 27721,
		437 => 27737,
		438 => 27754,
		439 => 27771,
		440 => 27787,
		441 => 27804,
		442 => 27820,
		443 => 27836,
		444 => 27853,
		445 => 27869,
		446 => 27885,
		447 => 27902,
		448 => 27918,
		449 => 27934,
		450 => 27950,
		451 => 27966,
		452 => 27982,
		453 => 27998,
		454 => 28014,
		455 => 28030,
		456 => 28045,
		457 => 28061,
		458 => 28077,
		459 => 28093,
		460 => 28108,
		461 => 28124,
		462 => 28139,
		463 => 28155,
		464 => 28170,
		465 => 28186,
		466 => 28201,
		467 => 28216,
		468 => 28232,
		469 => 28247,
		470 => 28262,
		471 => 28277,
		472 => 28292,
		473 => 28308,
		474 => 28323,
		475 => 28338,
		476 => 28353,
		477 => 28367,
		478 => 28382,
		479 => 28397,
		480 => 28412,
		481 => 28427,
		482 => 28441,
		483 => 28456,
		484 => 28471,
		485 => 28485,
		486 => 28500,
		487 => 28514,
		488 => 28529,
		489 => 28543,
		490 => 28557,
		491 => 28572,
		492 => 28586,
		493 => 28600,
		494 => 28614,
		495 => 28628,
		496 => 28643,
		497 => 28657,
		498 => 28671,
		499 => 28685,
		500 => 28699,
		501 => 28713,
		502 => 28726,
		503 => 28740,
		504 => 28754,
		505 => 28768,
		506 => 28781,
		507 => 28795,
		508 => 28809,
		509 => 28822,
		510 => 28836,
		511 => 28849,
		512 => 28863,
		513 => 28876,
		514 => 28890,
		515 => 28903,
		516 => 28916,
		517 => 28929,
		518 => 28943,
		519 => 28956,
		520 => 28969,
		521 => 28982,
		522 => 28995,
		523 => 29008,
		524 => 29021,
		525 => 29034,
		526 => 29047,
		527 => 29060,
		528 => 29073,
		529 => 29085,
		530 => 29098,
		531 => 29111,
		532 => 29124,
		533 => 29136,
		534 => 29149,
		535 => 29161,
		536 => 29174,
		537 => 29186,
		538 => 29199,
		539 => 29211,
		540 => 29224,
		541 => 29236,
		542 => 29248,
		543 => 29260,
		544 => 29273,
		545 => 29285,
		546 => 29297,
		547 => 29309,
		548 => 29321,
		549 => 29333,
		550 => 29345,
		551 => 29357,
		552 => 29369,
		553 => 29381,
		554 => 29393,
		555 => 29405,
		556 => 29416,
		557 => 29428,
		558 => 29440,
		559 => 29451,
		560 => 29463,
		561 => 29475,
		562 => 29486,
		563 => 29498,
		564 => 29509,
		565 => 29521,
		566 => 29532,
		567 => 29543,
		568 => 29555,
		569 => 29566,
		570 => 29577,
		571 => 29589,
		572 => 29600,
		573 => 29611,
		574 => 29622,
		575 => 29633,
		576 => 29644,
		577 => 29655,
		578 => 29666,
		579 => 29677,
		580 => 29688,
		581 => 29699,
		582 => 29710,
		583 => 29721,
		584 => 29731,
		585 => 29742,
		586 => 29753,
		587 => 29764,
		588 => 29774,
		589 => 29785,
		590 => 29795,
		591 => 29806,
		592 => 29816,
		593 => 29827,
		594 => 29837,
		595 => 29848,
		596 => 29858,
		597 => 29868,
		598 => 29879,
		599 => 29889,
		600 => 29899,
		601 => 29910,
		602 => 29920,
		603 => 29930,
		604 => 29940,
		605 => 29950,
		606 => 29960,
		607 => 29970,
		608 => 29980,
		609 => 29990,
		610 => 30000,
		611 => 30010,
		612 => 30020,
		613 => 30029,
		614 => 30039,
		615 => 30049,
		616 => 30059,
		617 => 30068,
		618 => 30078,
		619 => 30088,
		620 => 30097,
		621 => 30107,
		622 => 30116,
		623 => 30126,
		624 => 30135,
		625 => 30145,
		626 => 30154,
		627 => 30164,
		628 => 30173,
		629 => 30182,
		630 => 30192,
		631 => 30201,
		632 => 30210,
		633 => 30219,
		634 => 30228,
		635 => 30238,
		636 => 30247,
		637 => 30256,
		638 => 30265,
		639 => 30274,
		640 => 30283,
		641 => 30292,
		642 => 30301,
		643 => 30310,
		644 => 30318,
		645 => 30327,
		646 => 30336,
		647 => 30345,
		648 => 30354,
		649 => 30362,
		650 => 30371,
		651 => 30380,
		652 => 30388,
		653 => 30397,
		654 => 30405,
		655 => 30414,
		656 => 30423,
		657 => 30431,
		658 => 30439,
		659 => 30448,
		660 => 30456,
		661 => 30465,
		662 => 30473,
		663 => 30481,
		664 => 30490,
		665 => 30498,
		666 => 30506,
		667 => 30514,
		668 => 30523,
		669 => 30531,
		670 => 30539,
		671 => 30547,
		672 => 30555,
		673 => 30563,
		674 => 30571,
		675 => 30579,
		676 => 30587,
		677 => 30595,
		678 => 30603,
		679 => 30611,
		680 => 30619,
		681 => 30626,
		682 => 30634,
		683 => 30642,
		684 => 30650,
		685 => 30658,
		686 => 30665,
		687 => 30673,
		688 => 30681,
		689 => 30688,
		690 => 30696,
		691 => 30703,
		692 => 30711,
		693 => 30718,
		694 => 30726,
		695 => 30733,
		696 => 30741,
		697 => 30748,
		698 => 30756,
		699 => 30763,
		700 => 30770,
		701 => 30778,
		702 => 30785,
		703 => 30792,
		704 => 30799,
		705 => 30807,
		706 => 30814,
		707 => 30821,
		708 => 30828,
		709 => 30835,
		710 => 30842,
		711 => 30849,
		712 => 30856,
		713 => 30863,
		714 => 30870,
		715 => 30877,
		716 => 30884,
		717 => 30891,
		718 => 30898,
		719 => 30905,
		720 => 30912,
		721 => 30919,
		722 => 30926,
		723 => 30932,
		724 => 30939,
		725 => 30946,
		726 => 30952,
		727 => 30959,
		728 => 30966,
		729 => 30972,
		730 => 30979,
		731 => 30986,
		732 => 30992,
		733 => 30999,
		734 => 31005,
		735 => 31012,
		736 => 31018,
		737 => 31025,
		738 => 31031,
		739 => 31038,
		740 => 31044,
		741 => 31050,
		742 => 31057,
		743 => 31063,
		744 => 31069,
		745 => 31076,
		746 => 31082,
		747 => 31088,
		748 => 31094,
		749 => 31100,
		750 => 31107,
		751 => 31113,
		752 => 31119,
		753 => 31125,
		754 => 31131,
		755 => 31137,
		756 => 31143,
		757 => 31149,
		758 => 31155,
		759 => 31161,
		760 => 31167,
		761 => 31173,
		762 => 31179,
		763 => 31185,
		764 => 31191,
		765 => 31197,
		766 => 31202,
		767 => 31208,
		768 => 31214,
		769 => 31220,
		770 => 31226,
		771 => 31231,
		772 => 31237,
		773 => 31243,
		774 => 31248,
		775 => 31254,
		776 => 31260,
		777 => 31265,
		778 => 31271,
		779 => 31276,
		780 => 31282,
		781 => 31288,
		782 => 31293,
		783 => 31299,
		784 => 31304,
		785 => 31309,
		786 => 31315,
		787 => 31320,
		788 => 31326,
		789 => 31331,
		790 => 31336,
		791 => 31342,
		792 => 31347,
		793 => 31352,
		794 => 31358,
		795 => 31363,
		796 => 31368,
		797 => 31373,
		798 => 31379,
		799 => 31384,
		800 => 31389,
		801 => 31394,
		802 => 31399,
		803 => 31404,
		804 => 31409,
		805 => 31414,
		806 => 31420,
		807 => 31425,
		808 => 31430,
		809 => 31435,
		810 => 31440,
		811 => 31445,
		812 => 31450,
		813 => 31454,
		814 => 31459,
		815 => 31464,
		816 => 31469,
		817 => 31474,
		818 => 31479,
		819 => 31484,
		820 => 31488,
		821 => 31493,
		822 => 31498,
		823 => 31503,
		824 => 31508,
		825 => 31512,
		826 => 31517,
		827 => 31522,
		828 => 31526,
		829 => 31531,
		830 => 31536,
		831 => 31540,
		832 => 31545,
		833 => 31549,
		834 => 31554,
		835 => 31559,
		836 => 31563,
		837 => 31568,
		838 => 31572,
		839 => 31577,
		840 => 31581,
		841 => 31586,
		842 => 31590,
		843 => 31594,
		844 => 31599,
		845 => 31603,
		846 => 31608,
		847 => 31612,
		848 => 31616,
		849 => 31621,
		850 => 31625,
		851 => 31629,
		852 => 31634,
		853 => 31638,
		854 => 31642,
		855 => 31646,
		856 => 31651,
		857 => 31655,
		858 => 31659,
		859 => 31663,
		860 => 31667,
		861 => 31671,
		862 => 31676,
		863 => 31680,
		864 => 31684,
		865 => 31688,
		866 => 31692,
		867 => 31696,
		868 => 31700,
		869 => 31704,
		870 => 31708,
		871 => 31712,
		872 => 31716,
		873 => 31720,
		874 => 31724,
		875 => 31728,
		876 => 31732,
		877 => 31736,
		878 => 31740,
		879 => 31743,
		880 => 31747,
		881 => 31751,
		882 => 31755,
		883 => 31759,
		884 => 31763,
		885 => 31766,
		886 => 31770,
		887 => 31774,
		888 => 31778,
		889 => 31782,
		890 => 31785,
		891 => 31789,
		892 => 31793,
		893 => 31796,
		894 => 31800,
		895 => 31804,
		896 => 31807,
		897 => 31811,
		898 => 31815,
		899 => 31818,
		900 => 31822,
		901 => 31825,
		902 => 31829,
		903 => 31832,
		904 => 31836,
		905 => 31840,
		906 => 31843,
		907 => 31847,
		908 => 31850,
		909 => 31854,
		910 => 31857,
		911 => 31860,
		912 => 31864,
		913 => 31867,
		914 => 31871,
		915 => 31874,
		916 => 31878,
		917 => 31881,
		918 => 31884,
		919 => 31888,
		920 => 31891,
		921 => 31894,
		922 => 31898,
		923 => 31901,
		924 => 31904,
		925 => 31907,
		926 => 31911,
		927 => 31914,
		928 => 31917,
		929 => 31920,
		930 => 31924,
		931 => 31927,
		932 => 31930,
		933 => 31933,
		934 => 31936,
		935 => 31940,
		936 => 31943,
		937 => 31946,
		938 => 31949,
		939 => 31952,
		940 => 31955,
		941 => 31958,
		942 => 31961,
		943 => 31964,
		944 => 31967,
		945 => 31970,
		946 => 31974,
		947 => 31977,
		948 => 31980,
		949 => 31983,
		950 => 31986,
		951 => 31988,
		952 => 31991,
		953 => 31994,
		954 => 31997,
		955 => 32000,
		956 => 32003,
		957 => 32006,
		958 => 32009,
		959 => 32012,
		960 => 32015,
		961 => 32018,
		962 => 32020,
		963 => 32023,
		964 => 32026,
		965 => 32029,
		966 => 32032,
		967 => 32035,
		968 => 32037,
		969 => 32040,
		970 => 32043,
		971 => 32046,
		972 => 32048,
		973 => 32051,
		974 => 32054,
		975 => 32057,
		976 => 32059,
		977 => 32062,
		978 => 32065,
		979 => 32067,
		980 => 32070,
		981 => 32073,
		982 => 32075,
		983 => 32078,
		984 => 32081,
		985 => 32083,
		986 => 32086,
		987 => 32089,
		988 => 32091,
		989 => 32094,
		990 => 32096,
		991 => 32099,
		992 => 32101,
		993 => 32104,
		994 => 32106,
		995 => 32109,
		996 => 32112,
		997 => 32114,
		998 => 32117,
		999 => 32119,
		1000 => 32121,
		1001 => 32124,
		1002 => 32126,
		1003 => 32129,
		1004 => 32131,
		1005 => 32134,
		1006 => 32136,
		1007 => 32139,
		1008 => 32141,
		1009 => 32143,
		1010 => 32146,
		1011 => 32148,
		1012 => 32150,
		1013 => 32153,
		1014 => 32155,
		1015 => 32158,
		1016 => 32160,
		1017 => 32162,
		1018 => 32165,
		1019 => 32167,
		1020 => 32169,
		1021 => 32171,
		1022 => 32174,
		1023 => 32176,
		1024 => 32178,
		1025 => 32180,
		1026 => 32183,
		1027 => 32185,
		1028 => 32187,
		1029 => 32189,
		1030 => 32192,
		1031 => 32194,
		1032 => 32196,
		1033 => 32198,
		1034 => 32200,
		1035 => 32203,
		1036 => 32205,
		1037 => 32207,
		1038 => 32209,
		1039 => 32211,
		1040 => 32213,
		1041 => 32215,
		1042 => 32218,
		1043 => 32220,
		1044 => 32222,
		1045 => 32224,
		1046 => 32226,
		1047 => 32228,
		1048 => 32230,
		1049 => 32232,
		1050 => 32234,
		1051 => 32236,
		1052 => 32238,
		1053 => 32240,
		1054 => 32242,
		1055 => 32244,
		1056 => 32246,
		1057 => 32248,
		1058 => 32250,
		1059 => 32252,
		1060 => 32254,
		1061 => 32256,
		1062 => 32258,
		1063 => 32260,
		1064 => 32262,
		1065 => 32264,
		1066 => 32266,
		1067 => 32268,
		1068 => 32270,
		1069 => 32272,
		1070 => 32274,
		1071 => 32276,
		1072 => 32277,
		1073 => 32279,
		1074 => 32281,
		1075 => 32283,
		1076 => 32285,
		1077 => 32287,
		1078 => 32289,
		1079 => 32290,
		1080 => 32292,
		1081 => 32294,
		1082 => 32296,
		1083 => 32298,
		1084 => 32300,
		1085 => 32301,
		1086 => 32303,
		1087 => 32305,
		1088 => 32307,
		1089 => 32308,
		1090 => 32310,
		1091 => 32312,
		1092 => 32314,
		1093 => 32315,
		1094 => 32317,
		1095 => 32319,
		1096 => 32321,
		1097 => 32322,
		1098 => 32324,
		1099 => 32326,
		1100 => 32327,
		1101 => 32329,
		1102 => 32331,
		1103 => 32333,
		1104 => 32334,
		1105 => 32336,
		1106 => 32338,
		1107 => 32339,
		1108 => 32341,
		1109 => 32342,
		1110 => 32344,
		1111 => 32346,
		1112 => 32347,
		1113 => 32349,
		1114 => 32351,
		1115 => 32352,
		1116 => 32354,
		1117 => 32355,
		1118 => 32357,
		1119 => 32359,
		1120 => 32360,
		1121 => 32362,
		1122 => 32363,
		1123 => 32365,
		1124 => 32366,
		1125 => 32368,
		1126 => 32369,
		1127 => 32371,
		1128 => 32372,
		1129 => 32374,
		1130 => 32375,
		1131 => 32377,
		1132 => 32378,
		1133 => 32380,
		1134 => 32381,
		1135 => 32383,
		1136 => 32384,
		1137 => 32386,
		1138 => 32387,
		1139 => 32389,
		1140 => 32390,
		1141 => 32392,
		1142 => 32393,
		1143 => 32395,
		1144 => 32396,
		1145 => 32398,
		1146 => 32399,
		1147 => 32400,
		1148 => 32402,
		1149 => 32403,
		1150 => 32405,
		1151 => 32406,
		1152 => 32407,
		1153 => 32409,
		1154 => 32410,
		1155 => 32412,
		1156 => 32413,
		1157 => 32414,
		1158 => 32416,
		1159 => 32417,
		1160 => 32418,
		1161 => 32420,
		1162 => 32421,
		1163 => 32422,
		1164 => 32424,
		1165 => 32425,
		1166 => 32426,
		1167 => 32428,
		1168 => 32429,
		1169 => 32430,
		1170 => 32432,
		1171 => 32433,
		1172 => 32434,
		1173 => 32435,
		1174 => 32437,
		1175 => 32438,
		1176 => 32439,
		1177 => 32441,
		1178 => 32442,
		1179 => 32443,
		1180 => 32444,
		1181 => 32446,
		1182 => 32447,
		1183 => 32448,
		1184 => 32449,
		1185 => 32450,
		1186 => 32452,
		1187 => 32453,
		1188 => 32454,
		1189 => 32455,
		1190 => 32457,
		1191 => 32458,
		1192 => 32459,
		1193 => 32460,
		1194 => 32461,
		1195 => 32462,
		1196 => 32464,
		1197 => 32465,
		1198 => 32466,
		1199 => 32467,
		1200 => 32468,
		1201 => 32469,
		1202 => 32471,
		1203 => 32472,
		1204 => 32473,
		1205 => 32474,
		1206 => 32475,
		1207 => 32476,
		1208 => 32477,
		1209 => 32479,
		1210 => 32480,
		1211 => 32481,
		1212 => 32482,
		1213 => 32483,
		1214 => 32484,
		1215 => 32485,
		1216 => 32486,
		1217 => 32487,
		1218 => 32488,
		1219 => 32490,
		1220 => 32491,
		1221 => 32492,
		1222 => 32493,
		1223 => 32494,
		1224 => 32495,
		1225 => 32496,
		1226 => 32497,
		1227 => 32498,
		1228 => 32499,
		1229 => 32500,
		1230 => 32501,
		1231 => 32502,
		1232 => 32503,
		1233 => 32504,
		1234 => 32505,
		1235 => 32506,
		1236 => 32507,
		1237 => 32508,
		1238 => 32509,
		1239 => 32510,
		1240 => 32511,
		1241 => 32512,
		1242 => 32513,
		1243 => 32514,
		1244 => 32515,
		1245 => 32516,
		1246 => 32517,
		1247 => 32518,
		1248 => 32519,
		1249 => 32520,
		1250 => 32521,
		1251 => 32522,
		1252 => 32523,
		1253 => 32524,
		1254 => 32525,
		1255 => 32526,
		1256 => 32527,
		1257 => 32528,
		1258 => 32528,
		1259 => 32529,
		1260 => 32530,
		1261 => 32531,
		1262 => 32532,
		1263 => 32533,
		1264 => 32534,
		1265 => 32535,
		1266 => 32536,
		1267 => 32537,
		1268 => 32538,
		1269 => 32538,
		1270 => 32539,
		1271 => 32540,
		1272 => 32541,
		1273 => 32542,
		1274 => 32543,
		1275 => 32544,
		1276 => 32545,
		1277 => 32545,
		1278 => 32546,
		1279 => 32547,
		1280 => 32548,
		1281 => 32549,
		1282 => 32550,
		1283 => 32550,
		1284 => 32551,
		1285 => 32552,
		1286 => 32553,
		1287 => 32554,
		1288 => 32555,
		1289 => 32555,
		1290 => 32556,
		1291 => 32557,
		1292 => 32558,
		1293 => 32559,
		1294 => 32560,
		1295 => 32560,
		1296 => 32561,
		1297 => 32562,
		1298 => 32563,
		1299 => 32564,
		1300 => 32564,
		1301 => 32565,
		1302 => 32566,
		1303 => 32567,
		1304 => 32567,
		1305 => 32568,
		1306 => 32569,
		1307 => 32570,
		1308 => 32571,
		1309 => 32571,
		1310 => 32572,
		1311 => 32573,
		1312 => 32574,
		1313 => 32574,
		1314 => 32575,
		1315 => 32576,
		1316 => 32577,
		1317 => 32577,
		1318 => 32578,
		1319 => 32579,
		1320 => 32579,
		1321 => 32580,
		1322 => 32581,
		1323 => 32582,
		1324 => 32582,
		1325 => 32583,
		1326 => 32584,
		1327 => 32585,
		1328 => 32585,
		1329 => 32586,
		1330 => 32587,
		1331 => 32587,
		1332 => 32588,
		1333 => 32589,
		1334 => 32589,
		1335 => 32590,
		1336 => 32591,
		1337 => 32591,
		1338 => 32592,
		1339 => 32593,
		1340 => 32593,
		1341 => 32594,
		1342 => 32595,
		1343 => 32596,
		1344 => 32596,
		1345 => 32597,
		1346 => 32597,
		1347 => 32598,
		1348 => 32599,
		1349 => 32599,
		1350 => 32600,
		1351 => 32601,
		1352 => 32601,
		1353 => 32602,
		1354 => 32603,
		1355 => 32603,
		1356 => 32604,
		1357 => 32605,
		1358 => 32605,
		1359 => 32606,
		1360 => 32606,
		1361 => 32607,
		1362 => 32608,
		1363 => 32608,
		1364 => 32609,
		1365 => 32610,
		1366 => 32610,
		1367 => 32611,
		1368 => 32611,
		1369 => 32612,
		1370 => 32613,
		1371 => 32613,
		1372 => 32614,
		1373 => 32614,
		1374 => 32615,
		1375 => 32616,
		1376 => 32616,
		1377 => 32617,
		1378 => 32617,
		1379 => 32618,
		1380 => 32618,
		1381 => 32619,
		1382 => 32620,
		1383 => 32620,
		1384 => 32621,
		1385 => 32621,
		1386 => 32622,
		1387 => 32622,
		1388 => 32623,
		1389 => 32624,
		1390 => 32624,
		1391 => 32625,
		1392 => 32625,
		1393 => 32626,
		1394 => 32626,
		1395 => 32627,
		1396 => 32627,
		1397 => 32628,
		1398 => 32629,
		1399 => 32629,
		1400 => 32630,
		1401 => 32630,
		1402 => 32631,
		1403 => 32631,
		1404 => 32632,
		1405 => 32632,
		1406 => 32633,
		1407 => 32633,
		1408 => 32634,
		1409 => 32634,
		1410 => 32635,
		1411 => 32635,
		1412 => 32636,
		1413 => 32636,
		1414 => 32637,
		1415 => 32637,
		1416 => 32638,
		1417 => 32638,
		1418 => 32639,
		1419 => 32639,
		1420 => 32640,
		1421 => 32640,
		1422 => 32641,
		1423 => 32641,
		1424 => 32642,
		1425 => 32642,
		1426 => 32643,
		1427 => 32643,
		1428 => 32644,
		1429 => 32644,
		1430 => 32645,
		1431 => 32645,
		1432 => 32646,
		1433 => 32646,
		1434 => 32647,
		1435 => 32647,
		1436 => 32648,
		1437 => 32648,
		1438 => 32648,
		1439 => 32649,
		1440 => 32649,
		1441 => 32650,
		1442 => 32650,
		1443 => 32651,
		1444 => 32651,
		1445 => 32652,
		1446 => 32652,
		1447 => 32653,
		1448 => 32653,
		1449 => 32653,
		1450 => 32654,
		1451 => 32654,
		1452 => 32655,
		1453 => 32655,
		1454 => 32656,
		1455 => 32656,
		1456 => 32657,
		1457 => 32657,
		1458 => 32657,
		1459 => 32658,
		1460 => 32658,
		1461 => 32659,
		1462 => 32659,
		1463 => 32659,
		1464 => 32660,
		1465 => 32660,
		1466 => 32661,
		1467 => 32661,
		1468 => 32662,
		1469 => 32662,
		1470 => 32662,
		1471 => 32663,
		1472 => 32663,
		1473 => 32664,
		1474 => 32664,
		1475 => 32664,
		1476 => 32665,
		1477 => 32665,
		1478 => 32666,
		1479 => 32666,
		1480 => 32666,
		1481 => 32667,
		1482 => 32667,
		1483 => 32668,
		1484 => 32668,
		1485 => 32668,
		1486 => 32669,
		1487 => 32669,
		1488 => 32669,
		1489 => 32670,
		1490 => 32670,
		1491 => 32671,
		1492 => 32671,
		1493 => 32671,
		1494 => 32672,
		1495 => 32672,
		1496 => 32672,
		1497 => 32673,
		1498 => 32673,
		1499 => 32674,
		1500 => 32674,
		1501 => 32674,
		1502 => 32675,
		1503 => 32675,
		1504 => 32675,
		1505 => 32676,
		1506 => 32676,
		1507 => 32676,
		1508 => 32677,
		1509 => 32677,
		1510 => 32677,
		1511 => 32678,
		1512 => 32678,
		1513 => 32679,
		1514 => 32679,
		1515 => 32679,
		1516 => 32680,
		1517 => 32680,
		1518 => 32680,
		1519 => 32681,
		1520 => 32681,
		1521 => 32681,
		1522 => 32682,
		1523 => 32682,
		1524 => 32682,
		1525 => 32683,
		1526 => 32683,
		1527 => 32683,
		1528 => 32684,
		1529 => 32684,
		1530 => 32684,
		1531 => 32685,
		1532 => 32685,
		1533 => 32685,
		1534 => 32685,
		1535 => 32686,
		1536 => 32686,
		1537 => 32686,
		1538 => 32687,
		1539 => 32687,
		1540 => 32687,
		1541 => 32688,
		1542 => 32688,
		1543 => 32688,
		1544 => 32689,
		1545 => 32689,
		1546 => 32689,
		1547 => 32689,
		1548 => 32690,
		1549 => 32690,
		1550 => 32690,
		1551 => 32691,
		1552 => 32691,
		1553 => 32691,
		1554 => 32692,
		1555 => 32692,
		1556 => 32692,
		1557 => 32692,
		1558 => 32693,
		1559 => 32693,
		1560 => 32693,
		1561 => 32694,
		1562 => 32694,
		1563 => 32694,
		1564 => 32694,
		1565 => 32695,
		1566 => 32695,
		1567 => 32695,
		1568 => 32696,
		1569 => 32696,
		1570 => 32696,
		1571 => 32696,
		1572 => 32697,
		1573 => 32697,
		1574 => 32697,
		1575 => 32698,
		1576 => 32698,
		1577 => 32698,
		1578 => 32698,
		1579 => 32699,
		1580 => 32699,
		1581 => 32699,
		1582 => 32699,
		1583 => 32700,
		1584 => 32700,
		1585 => 32700,
		1586 => 32700,
		1587 => 32701,
		1588 => 32701,
		1589 => 32701,
		1590 => 32701,
		1591 => 32702,
		1592 => 32702,
		1593 => 32702,
		1594 => 32702,
		1595 => 32703,
		1596 => 32703,
		1597 => 32703,
		1598 => 32703,
		1599 => 32704,
		1600 => 32704,
		1601 => 32704,
		1602 => 32704,
		1603 => 32705,
		1604 => 32705,
		1605 => 32705,
		1606 => 32705,
		1607 => 32706,
		1608 => 32706,
		1609 => 32706,
		1610 => 32706,
		1611 => 32707,
		1612 => 32707,
		1613 => 32707,
		1614 => 32707,
		1615 => 32708,
		1616 => 32708,
		1617 => 32708,
		1618 => 32708,
		1619 => 32708,
		1620 => 32709,
		1621 => 32709,
		1622 => 32709,
		1623 => 32709,
		1624 => 32710,
		1625 => 32710,
		1626 => 32710,
		1627 => 32710,
		1628 => 32710,
		1629 => 32711,
		1630 => 32711,
		1631 => 32711,
		1632 => 32711,
		1633 => 32712,
		1634 => 32712,
		1635 => 32712,
		1636 => 32712,
		1637 => 32712,
		1638 => 32713,
		1639 => 32713,
		1640 => 32713,
		1641 => 32713,
		1642 => 32713,
		1643 => 32714,
		1644 => 32714,
		1645 => 32714,
		1646 => 32714,
		1647 => 32715,
		1648 => 32715,
		1649 => 32715,
		1650 => 32715,
		1651 => 32715,
		1652 => 32716,
		1653 => 32716,
		1654 => 32716,
		1655 => 32716,
		1656 => 32716,
		1657 => 32717,
		1658 => 32717,
		1659 => 32717,
		1660 => 32717,
		1661 => 32717,
		1662 => 32718,
		1663 => 32718,
		1664 => 32718,
		1665 => 32718,
		1666 => 32718,
		1667 => 32718,
		1668 => 32719,
		1669 => 32719,
		1670 => 32719,
		1671 => 32719,
		1672 => 32719,
		1673 => 32720,
		1674 => 32720,
		1675 => 32720,
		1676 => 32720,
		1677 => 32720,
		1678 => 32720,
		1679 => 32721,
		1680 => 32721,
		1681 => 32721,
		1682 => 32721,
		1683 => 32721,
		1684 => 32722,
		1685 => 32722,
		1686 => 32722,
		1687 => 32722,
		1688 => 32722,
		1689 => 32722,
		1690 => 32723,
		1691 => 32723,
		1692 => 32723,
		1693 => 32723,
		1694 => 32723,
		1695 => 32723,
		1696 => 32724,
		1697 => 32724,
		1698 => 32724,
		1699 => 32724,
		1700 => 32724,
		1701 => 32724,
		1702 => 32725,
		1703 => 32725,
		1704 => 32725,
		1705 => 32725,
		1706 => 32725,
		1707 => 32725,
		1708 => 32726,
		1709 => 32726,
		1710 => 32726,
		1711 => 32726,
		1712 => 32726,
		1713 => 32726,
		1714 => 32727,
		1715 => 32727,
		1716 => 32727,
		1717 => 32727,
		1718 => 32727,
		1719 => 32727,
		1720 => 32728,
		1721 => 32728,
		1722 => 32728,
		1723 => 32728,
		1724 => 32728,
		1725 => 32728,
		1726 => 32728,
		1727 => 32729,
		1728 => 32729,
		1729 => 32729,
		1730 => 32729,
		1731 => 32729,
		1732 => 32729,
		1733 => 32729,
		1734 => 32730,
		1735 => 32730,
		1736 => 32730,
		1737 => 32730,
		1738 => 32730,
		1739 => 32730,
		1740 => 32730,
		1741 => 32731,
		1742 => 32731,
		1743 => 32731,
		1744 => 32731,
		1745 => 32731,
		1746 => 32731,
		1747 => 32731,
		1748 => 32732,
		1749 => 32732,
		1750 => 32732,
		1751 => 32732,
		1752 => 32732,
		1753 => 32732,
		1754 => 32732,
		1755 => 32733,
		1756 => 32733,
		1757 => 32733,
		1758 => 32733,
		1759 => 32733,
		1760 => 32733,
		1761 => 32733,
		1762 => 32733,
		1763 => 32734,
		1764 => 32734,
		1765 => 32734,
		1766 => 32734,
		1767 => 32734,
		1768 => 32734,
		1769 => 32734,
		1770 => 32735,
		1771 => 32735,
		1772 => 32735,
		1773 => 32735,
		1774 => 32735,
		1775 => 32735,
		1776 => 32735,
		1777 => 32735,
		1778 => 32736,
		1779 => 32736,
		1780 => 32736,
		1781 => 32736,
		1782 => 32736,
		1783 => 32736,
		1784 => 32736,
		1785 => 32736,
		1786 => 32736,
		1787 => 32737,
		1788 => 32737,
		1789 => 32737,
		1790 => 32737,
		1791 => 32737,
		1792 => 32737,
		1793 => 32737,
		1794 => 32737,
		1795 => 32738,
		1796 => 32738,
		1797 => 32738,
		1798 => 32738,
		1799 => 32738,
		1800 => 32738,
		1801 => 32738,
		1802 => 32738,
		1803 => 32738,
		1804 => 32739,
		1805 => 32739,
		1806 => 32739,
		1807 => 32739,
		1808 => 32739,
		1809 => 32739,
		1810 => 32739,
		1811 => 32739,
		1812 => 32739,
		1813 => 32740,
		1814 => 32740,
		1815 => 32740,
		1816 => 32740,
		1817 => 32740,
		1818 => 32740,
		1819 => 32740,
		1820 => 32740,
		1821 => 32740,
		1822 => 32740,
		1823 => 32741,
		1824 => 32741,
		1825 => 32741,
		1826 => 32741,
		1827 => 32741,
		1828 => 32741,
		1829 => 32741,
		1830 => 32741,
		1831 => 32741,
		1832 => 32742,
		1833 => 32742,
		1834 => 32742,
		1835 => 32742,
		1836 => 32742,
		1837 => 32742,
		1838 => 32742,
		1839 => 32742,
		1840 => 32742,
		1841 => 32742,
		1842 => 32742,
		1843 => 32743,
		1844 => 32743,
		1845 => 32743,
		1846 => 32743,
		1847 => 32743,
		1848 => 32743,
		1849 => 32743,
		1850 => 32743,
		1851 => 32743,
		1852 => 32743,
		1853 => 32744,
		1854 => 32744,
		1855 => 32744,
		1856 => 32744,
		1857 => 32744,
		1858 => 32744,
		1859 => 32744,
		1860 => 32744,
		1861 => 32744,
		1862 => 32744,
		1863 => 32744,
		1864 => 32745,
		1865 => 32745,
		1866 => 32745,
		1867 => 32745,
		1868 => 32745,
		1869 => 32745,
		1870 => 32745,
		1871 => 32745,
		1872 => 32745,
		1873 => 32745,
		1874 => 32745,
		1875 => 32745,
		1876 => 32746,
		1877 => 32746,
		1878 => 32746,
		1879 => 32746,
		1880 => 32746,
		1881 => 32746,
		1882 => 32746,
		1883 => 32746,
		1884 => 32746,
		1885 => 32746,
		1886 => 32746,
		1887 => 32746,
		1888 => 32747,
		1889 => 32747,
		1890 => 32747,
		1891 => 32747,
		1892 => 32747,
		1893 => 32747,
		1894 => 32747,
		1895 => 32747,
		1896 => 32747,
		1897 => 32747,
		1898 => 32747,
		1899 => 32747,
		1900 => 32747,
		1901 => 32748,
		1902 => 32748,
		1903 => 32748,
		1904 => 32748,
		1905 => 32748,
		1906 => 32748,
		1907 => 32748,
		1908 => 32748,
		1909 => 32748,
		1910 => 32748,
		1911 => 32748,
		1912 => 32748,
		1913 => 32748,
		1914 => 32748,
		1915 => 32749,
		1916 => 32749,
		1917 => 32749,
		1918 => 32749,
		1919 => 32749,
		1920 => 32749,
		1921 => 32749,
		1922 => 32749,
		1923 => 32749,
		1924 => 32749,
		1925 => 32749,
		1926 => 32749,
		1927 => 32749,
		1928 => 32749,
		1929 => 32750,
		1930 => 32750,
		1931 => 32750,
		1932 => 32750,
		1933 => 32750,
		1934 => 32750,
		1935 => 32750,
		1936 => 32750,
		1937 => 32750,
		1938 => 32750,
		1939 => 32750,
		1940 => 32750,
		1941 => 32750,
		1942 => 32750,
		1943 => 32750,
		1944 => 32751,
		1945 => 32751,
		1946 => 32751,
		1947 => 32751,
		1948 => 32751,
		1949 => 32751,
		1950 => 32751,
		1951 => 32751,
		1952 => 32751,
		1953 => 32751,
		1954 => 32751,
		1955 => 32751,
		1956 => 32751,
		1957 => 32751,
		1958 => 32751,
		1959 => 32751,
		1960 => 32752,
		1961 => 32752,
		1962 => 32752,
		1963 => 32752,
		1964 => 32752,
		1965 => 32752,
		1966 => 32752,
		1967 => 32752,
		1968 => 32752,
		1969 => 32752,
		1970 => 32752,
		1971 => 32752,
		1972 => 32752,
		1973 => 32752,
		1974 => 32752,
		1975 => 32752,
		1976 => 32752,
		1977 => 32753,
		1978 => 32753,
		1979 => 32753,
		1980 => 32753,
		1981 => 32753,
		1982 => 32753,
		1983 => 32753,
		1984 => 32753,
		1985 => 32753,
		1986 => 32753,
		1987 => 32753,
		1988 => 32753,
		1989 => 32753,
		1990 => 32753,
		1991 => 32753,
		1992 => 32753,
		1993 => 32753,
		1994 => 32753,
		1995 => 32754,
		1996 => 32754,
		1997 => 32754,
		1998 => 32754,
		1999 => 32754,
		2000 => 32754,
		2001 => 32754,
		2002 => 32754,
		2003 => 32754,
		2004 => 32754,
		2005 => 32754,
		2006 => 32754,
		2007 => 32754,
		2008 => 32754,
		2009 => 32754,
		2010 => 32754,
		2011 => 32754,
		2012 => 32754,
		2013 => 32754,
		2014 => 32754,
		2015 => 32755,
		2016 => 32755,
		2017 => 32755,
		2018 => 32755,
		2019 => 32755,
		2020 => 32755,
		2021 => 32755,
		2022 => 32755,
		2023 => 32755,
		2024 => 32755,
		2025 => 32755,
		2026 => 32755,
		2027 => 32755,
		2028 => 32755,
		2029 => 32755,
		2030 => 32755,
		2031 => 32755,
		2032 => 32755,
		2033 => 32755,
		2034 => 32755,
		2035 => 32755,
		2036 => 32756,
		2037 => 32756,
		2038 => 32756,
		2039 => 32756,
		2040 => 32756,
		2041 => 32756,
		2042 => 32756,
		2043 => 32756,
		2044 => 32756,
		2045 => 32756,
		2046 => 32756,
		2047 => 32756,
		2048 => 32756,
		2049 => 32756,
		2050 => 32756,
		2051 => 32756,
		2052 => 32756,
		2053 => 32756,
		2054 => 32756,
		2055 => 32756,
		2056 => 32756,
		2057 => 32756,
		2058 => 32756,
		2059 => 32756,
		2060 => 32757,
		2061 => 32757,
		2062 => 32757,
		2063 => 32757,
		2064 => 32757,
		2065 => 32757,
		2066 => 32757,
		2067 => 32757,
		2068 => 32757,
		2069 => 32757,
		2070 => 32757,
		2071 => 32757,
		2072 => 32757,
		2073 => 32757,
		2074 => 32757,
		2075 => 32757,
		2076 => 32757,
		2077 => 32757,
		2078 => 32757,
		2079 => 32757,
		2080 => 32757,
		2081 => 32757,
		2082 => 32757,
		2083 => 32757,
		2084 => 32757,
		2085 => 32758,
		2086 => 32758,
		2087 => 32758,
		2088 => 32758,
		2089 => 32758,
		2090 => 32758,
		2091 => 32758,
		2092 => 32758,
		2093 => 32758,
		2094 => 32758,
		2095 => 32758,
		2096 => 32758,
		2097 => 32758,
		2098 => 32758,
		2099 => 32758,
		2100 => 32758,
		2101 => 32758,
		2102 => 32758,
		2103 => 32758,
		2104 => 32758,
		2105 => 32758,
		2106 => 32758,
		2107 => 32758,
		2108 => 32758,
		2109 => 32758,
		2110 => 32758,
		2111 => 32758,
		2112 => 32758,
		2113 => 32758,
		2114 => 32759,
		2115 => 32759,
		2116 => 32759,
		2117 => 32759,
		2118 => 32759,
		2119 => 32759,
		2120 => 32759,
		2121 => 32759,
		2122 => 32759,
		2123 => 32759,
		2124 => 32759,
		2125 => 32759,
		2126 => 32759,
		2127 => 32759,
		2128 => 32759,
		2129 => 32759,
		2130 => 32759,
		2131 => 32759,
		2132 => 32759,
		2133 => 32759,
		2134 => 32759,
		2135 => 32759,
		2136 => 32759,
		2137 => 32759,
		2138 => 32759,
		2139 => 32759,
		2140 => 32759,
		2141 => 32759,
		2142 => 32759,
		2143 => 32759,
		2144 => 32759,
		2145 => 32759,
		2146 => 32760,
		2147 => 32760,
		2148 => 32760,
		2149 => 32760,
		2150 => 32760,
		2151 => 32760,
		2152 => 32760,
		2153 => 32760,
		2154 => 32760,
		2155 => 32760,
		2156 => 32760,
		2157 => 32760,
		2158 => 32760,
		2159 => 32760,
		2160 => 32760,
		2161 => 32760,
		2162 => 32760,
		2163 => 32760,
		2164 => 32760,
		2165 => 32760,
		2166 => 32760,
		2167 => 32760,
		2168 => 32760,
		2169 => 32760,
		2170 => 32760,
		2171 => 32760,
		2172 => 32760,
		2173 => 32760,
		2174 => 32760,
		2175 => 32760,
		2176 => 32760,
		2177 => 32760,
		2178 => 32760,
		2179 => 32760,
		2180 => 32760,
		2181 => 32760,
		2182 => 32761,
		2183 => 32761,
		2184 => 32761,
		2185 => 32761,
		2186 => 32761,
		2187 => 32761,
		2188 => 32761,
		2189 => 32761,
		2190 => 32761,
		2191 => 32761,
		2192 => 32761,
		2193 => 32761,
		2194 => 32761,
		2195 => 32761,
		2196 => 32761,
		2197 => 32761,
		2198 => 32761,
		2199 => 32761,
		2200 => 32761,
		2201 => 32761,
		2202 => 32761,
		2203 => 32761,
		2204 => 32761,
		2205 => 32761,
		2206 => 32761,
		2207 => 32761,
		2208 => 32761,
		2209 => 32761,
		2210 => 32761,
		2211 => 32761,
		2212 => 32761,
		2213 => 32761,
		2214 => 32761,
		2215 => 32761,
		2216 => 32761,
		2217 => 32761,
		2218 => 32761,
		2219 => 32761,
		2220 => 32761,
		2221 => 32761,
		2222 => 32761,
		2223 => 32761,
		2224 => 32761,
		2225 => 32762,
		2226 => 32762,
		2227 => 32762,
		2228 => 32762,
		2229 => 32762,
		2230 => 32762,
		2231 => 32762,
		2232 => 32762,
		2233 => 32762,
		2234 => 32762,
		2235 => 32762,
		2236 => 32762,
		2237 => 32762,
		2238 => 32762,
		2239 => 32762,
		2240 => 32762,
		2241 => 32762,
		2242 => 32762,
		2243 => 32762,
		2244 => 32762,
		2245 => 32762,
		2246 => 32762,
		2247 => 32762,
		2248 => 32762,
		2249 => 32762,
		2250 => 32762,
		2251 => 32762,
		2252 => 32762,
		2253 => 32762,
		2254 => 32762,
		2255 => 32762,
		2256 => 32762,
		2257 => 32762,
		2258 => 32762,
		2259 => 32762,
		2260 => 32762,
		2261 => 32762,
		2262 => 32762,
		2263 => 32762,
		2264 => 32762,
		2265 => 32762,
		2266 => 32762,
		2267 => 32762,
		2268 => 32762,
		2269 => 32762,
		2270 => 32762,
		2271 => 32762,
		2272 => 32762,
		2273 => 32762,
		2274 => 32762,
		2275 => 32762,
		2276 => 32762,
		2277 => 32763,
		2278 => 32763,
		2279 => 32763,
		2280 => 32763,
		2281 => 32763,
		2282 => 32763,
		2283 => 32763,
		2284 => 32763,
		2285 => 32763,
		2286 => 32763,
		2287 => 32763,
		2288 => 32763,
		2289 => 32763,
		2290 => 32763,
		2291 => 32763,
		2292 => 32763,
		2293 => 32763,
		2294 => 32763,
		2295 => 32763,
		2296 => 32763,
		2297 => 32763,
		2298 => 32763,
		2299 => 32763,
		2300 => 32763,
		2301 => 32763,
		2302 => 32763,
		2303 => 32763,
		2304 => 32763,
		2305 => 32763,
		2306 => 32763,
		2307 => 32763,
		2308 => 32763,
		2309 => 32763,
		2310 => 32763,
		2311 => 32763,
		2312 => 32763,
		2313 => 32763,
		2314 => 32763,
		2315 => 32763,
		2316 => 32763,
		2317 => 32763,
		2318 => 32763,
		2319 => 32763,
		2320 => 32763,
		2321 => 32763,
		2322 => 32763,
		2323 => 32763,
		2324 => 32763,
		2325 => 32763,
		2326 => 32763,
		2327 => 32763,
		2328 => 32763,
		2329 => 32763,
		2330 => 32763,
		2331 => 32763,
		2332 => 32763,
		2333 => 32763,
		2334 => 32763,
		2335 => 32763,
		2336 => 32763,
		2337 => 32763,
		2338 => 32763,
		2339 => 32763,
		2340 => 32763,
		2341 => 32764,
		2342 => 32764,
		2343 => 32764,
		2344 => 32764,
		2345 => 32764,
		2346 => 32764,
		2347 => 32764,
		2348 => 32764,
		2349 => 32764,
		2350 => 32764,
		2351 => 32764,
		2352 => 32764,
		2353 => 32764,
		2354 => 32764,
		2355 => 32764,
		2356 => 32764,
		2357 => 32764,
		2358 => 32764,
		2359 => 32764,
		2360 => 32764,
		2361 => 32764,
		2362 => 32764,
		2363 => 32764,
		2364 => 32764,
		2365 => 32764,
		2366 => 32764,
		2367 => 32764,
		2368 => 32764,
		2369 => 32764,
		2370 => 32764,
		2371 => 32764,
		2372 => 32764,
		2373 => 32764,
		2374 => 32764,
		2375 => 32764,
		2376 => 32764,
		2377 => 32764,
		2378 => 32764,
		2379 => 32764,
		2380 => 32764,
		2381 => 32764,
		2382 => 32764,
		2383 => 32764,
		2384 => 32764,
		2385 => 32764,
		2386 => 32764,
		2387 => 32764,
		2388 => 32764,
		2389 => 32764,
		2390 => 32764,
		2391 => 32764,
		2392 => 32764,
		2393 => 32764,
		2394 => 32764,
		2395 => 32764,
		2396 => 32764,
		2397 => 32764,
		2398 => 32764,
		2399 => 32764,
		2400 => 32764,
		2401 => 32764,
		2402 => 32764,
		2403 => 32764,
		2404 => 32764,
		2405 => 32764,
		2406 => 32764,
		2407 => 32764,
		2408 => 32764,
		2409 => 32764,
		2410 => 32764,
		2411 => 32764,
		2412 => 32764,
		2413 => 32764,
		2414 => 32764,
		2415 => 32764,
		2416 => 32764,
		2417 => 32764,
		2418 => 32764,
		2419 => 32764,
		2420 => 32764,
		2421 => 32764,
		2422 => 32764,
		2423 => 32764,
		2424 => 32764,
		2425 => 32764,
		2426 => 32764,
		2427 => 32765,
		2428 => 32765,
		2429 => 32765,
		2430 => 32765,
		2431 => 32765,
		2432 => 32765,
		2433 => 32765,
		2434 => 32765,
		2435 => 32765,
		2436 => 32765,
		2437 => 32765,
		2438 => 32765,
		2439 => 32765,
		2440 => 32765,
		2441 => 32765,
		2442 => 32765,
		2443 => 32765,
		2444 => 32765,
		2445 => 32765,
		2446 => 32765,
		2447 => 32765,
		2448 => 32765,
		2449 => 32765,
		2450 => 32765,
		2451 => 32765,
		2452 => 32765,
		2453 => 32765,
		2454 => 32765,
		2455 => 32765,
		2456 => 32765,
		2457 => 32765,
		2458 => 32765,
		2459 => 32765,
		2460 => 32765,
		2461 => 32765,
		2462 => 32765,
		2463 => 32765,
		2464 => 32765,
		2465 => 32765,
		2466 => 32765,
		2467 => 32765,
		2468 => 32765,
		2469 => 32765,
		2470 => 32765,
		2471 => 32765,
		2472 => 32765,
		2473 => 32765,
		2474 => 32765,
		2475 => 32765,
		2476 => 32765,
		2477 => 32765,
		2478 => 32765,
		2479 => 32765,
		2480 => 32765,
		2481 => 32765,
		2482 => 32765,
		2483 => 32765,
		2484 => 32765,
		2485 => 32765,
		2486 => 32765,
		2487 => 32765,
		2488 => 32765,
		2489 => 32765,
		2490 => 32765,
		2491 => 32765,
		2492 => 32765,
		2493 => 32765,
		2494 => 32765,
		2495 => 32765,
		2496 => 32765,
		2497 => 32765,
		2498 => 32765,
		2499 => 32765,
		2500 => 32765,
		2501 => 32765,
		2502 => 32765,
		2503 => 32765,
		2504 => 32765,
		2505 => 32765,
		2506 => 32765,
		2507 => 32765,
		2508 => 32765,
		2509 => 32765,
		2510 => 32765,
		2511 => 32765,
		2512 => 32765,
		2513 => 32765,
		2514 => 32765,
		2515 => 32765,
		2516 => 32765,
		2517 => 32765,
		2518 => 32765,
		2519 => 32765,
		2520 => 32765,
		2521 => 32765,
		2522 => 32765,
		2523 => 32765,
		2524 => 32765,
		2525 => 32765,
		2526 => 32765,
		2527 => 32765,
		2528 => 32765,
		2529 => 32765,
		2530 => 32765,
		2531 => 32765,
		2532 => 32765,
		2533 => 32765,
		2534 => 32765,
		2535 => 32765,
		2536 => 32765,
		2537 => 32765,
		2538 => 32765,
		2539 => 32765,
		2540 => 32765,
		2541 => 32765,
		2542 => 32765,
		2543 => 32765,
		2544 => 32765,
		2545 => 32765,
		2546 => 32765,
		2547 => 32765,
		2548 => 32765,
		2549 => 32765,
		2550 => 32765,
		2551 => 32765,
		2552 => 32765,
		2553 => 32765,
		2554 => 32765,
		2555 => 32765,
		2556 => 32765,
		2557 => 32765,
		2558 => 32766,
		2559 => 32766,
		2560 => 32766,
		2561 => 32766,
		2562 => 32766,
		2563 => 32766,
		2564 => 32766,
		2565 => 32766,
		2566 => 32766,
		2567 => 32766,
		2568 => 32766,
		2569 => 32766,
		2570 => 32766,
		2571 => 32766,
		2572 => 32766,
		2573 => 32766,
		2574 => 32766,
		2575 => 32766,
		2576 => 32766,
		2577 => 32766,
		2578 => 32766,
		2579 => 32766,
		2580 => 32766,
		2581 => 32766,
		2582 => 32766,
		2583 => 32766,
		2584 => 32766,
		2585 => 32766,
		2586 => 32766,
		2587 => 32766,
		2588 => 32766,
		2589 => 32766,
		2590 => 32766,
		2591 => 32766,
		2592 => 32766,
		2593 => 32766,
		2594 => 32766,
		2595 => 32766,
		2596 => 32766,
		2597 => 32766,
		2598 => 32766,
		2599 => 32766,
		2600 => 32766,
		2601 => 32766,
		2602 => 32766,
		2603 => 32766,
		2604 => 32766,
		2605 => 32766,
		2606 => 32766,
		2607 => 32766,
		2608 => 32766,
		2609 => 32766,
		2610 => 32766,
		2611 => 32766,
		2612 => 32766,
		2613 => 32766,
		2614 => 32766,
		2615 => 32766,
		2616 => 32766,
		2617 => 32766,
		2618 => 32766,
		2619 => 32766,
		2620 => 32766,
		2621 => 32766,
		2622 => 32766,
		2623 => 32766,
		2624 => 32766,
		2625 => 32766,
		2626 => 32766,
		2627 => 32766,
		2628 => 32766,
		2629 => 32766,
		2630 => 32766,
		2631 => 32766,
		2632 => 32766,
		2633 => 32766,
		2634 => 32766,
		2635 => 32766,
		2636 => 32766,
		2637 => 32766,
		2638 => 32766,
		2639 => 32766,
		2640 => 32766,
		2641 => 32766,
		2642 => 32766,
		2643 => 32766,
		2644 => 32766,
		2645 => 32766,
		2646 => 32766,
		2647 => 32766,
		2648 => 32766,
		2649 => 32766,
		2650 => 32766,
		2651 => 32766,
		2652 => 32766,
		2653 => 32766,
		2654 => 32766,
		2655 => 32766,
		2656 => 32766,
		2657 => 32766,
		2658 => 32766,
		2659 => 32766,
		2660 => 32766,
		2661 => 32766,
		2662 => 32766,
		2663 => 32766,
		2664 => 32766,
		2665 => 32766,
		2666 => 32766,
		2667 => 32766,
		2668 => 32766,
		2669 => 32766,
		2670 => 32766,
		2671 => 32766,
		2672 => 32766,
		2673 => 32766,
		2674 => 32766,
		2675 => 32766,
		2676 => 32766,
		2677 => 32766,
		2678 => 32766,
		2679 => 32766,
		2680 => 32766,
		2681 => 32766,
		2682 => 32766,
		2683 => 32766,
		2684 => 32766,
		2685 => 32766,
		2686 => 32766,
		2687 => 32766,
		2688 => 32766,
		2689 => 32766,
		2690 => 32766,
		2691 => 32766,
		2692 => 32766,
		2693 => 32766,
		2694 => 32766,
		2695 => 32766,
		2696 => 32766,
		2697 => 32766,
		2698 => 32766,
		2699 => 32766,
		2700 => 32766,
		2701 => 32766,
		2702 => 32766,
		2703 => 32766,
		2704 => 32766,
		2705 => 32766,
		2706 => 32766,
		2707 => 32766,
		2708 => 32766,
		2709 => 32766,
		2710 => 32766,
		2711 => 32766,
		2712 => 32766,
		2713 => 32766,
		2714 => 32766,
		2715 => 32766,
		2716 => 32766,
		2717 => 32766,
		2718 => 32766,
		2719 => 32766,
		2720 => 32766,
		2721 => 32766,
		2722 => 32766,
		2723 => 32766,
		2724 => 32766,
		2725 => 32766,
		2726 => 32766,
		2727 => 32766,
		2728 => 32766,
		2729 => 32766,
		2730 => 32766,
		2731 => 32766,
		2732 => 32766,
		2733 => 32766,
		2734 => 32766,
		2735 => 32766,
		2736 => 32766,
		2737 => 32766,
		2738 => 32766,
		2739 => 32766,
		2740 => 32766,
		2741 => 32766,
		2742 => 32766,
		2743 => 32766,
		2744 => 32766,
		2745 => 32766,
		2746 => 32766,
		2747 => 32766,
		2748 => 32766,
		2749 => 32766,
		2750 => 32766,
		2751 => 32766,
		2752 => 32766,
		2753 => 32766,
		2754 => 32766,
		2755 => 32766,
		2756 => 32766,
		2757 => 32766,
		2758 => 32766,
		2759 => 32766,
		2760 => 32766,
		2761 => 32766,
		2762 => 32766,
		2763 => 32766,
		2764 => 32766,
		2765 => 32766,
		2766 => 32766,
		2767 => 32766,
		2768 => 32766,
		2769 => 32766,
		2770 => 32766,
		2771 => 32766,
		2772 => 32766,
		2773 => 32766,
		2774 => 32766,
		2775 => 32766,
		2776 => 32766,
		2777 => 32766,
		2778 => 32766,
		2779 => 32766,
		2780 => 32766,
		2781 => 32766,
		2782 => 32766,
		2783 => 32766,
		2784 => 32766,
		2785 => 32766,
		2786 => 32766,
		2787 => 32766,
		2788 => 32766,
		2789 => 32766,
		2790 => 32766,
		2791 => 32766,
		2792 => 32766,
		2793 => 32766,
		2794 => 32766,
		2795 => 32766,
		2796 => 32766,
		2797 => 32766,
		2798 => 32766,
		2799 => 32766,
		2800 => 32766,
		2801 => 32766,
		2802 => 32766,
		2803 => 32766,
		2804 => 32766,
		2805 => 32766,
		2806 => 32766,
		2807 => 32766,
		2808 => 32766,
		2809 => 32766,
		2810 => 32766,
		2811 => 32766,
		2812 => 32766,
		2813 => 32766,
		2814 => 32766,
		2815 => 32766,
		2816 => 32766,
		2817 => 32766,
		2818 => 32766,
		2819 => 32766,
		2820 => 32766,
		2821 => 32766,
		2822 => 32766,
		2823 => 32766,
		2824 => 32766,
		2825 => 32766,
		2826 => 32766,
		2827 => 32766,
		2828 => 32766,
		2829 => 32766,
		2830 => 32766,
		2831 => 32766,
		2832 => 32766,
		2833 => 32766,
		2834 => 32766,
		2835 => 32766,
		2836 => 32766,
		2837 => 32766,
		2838 => 32766,
		2839 => 32767,
		2840 => 32767,
		2841 => 32767,
		2842 => 32767,
		2843 => 32767,
		2844 => 32767,
		2845 => 32767,
		2846 => 32767,
		2847 => 32767,
		2848 => 32767,
		2849 => 32767,
		2850 => 32767,
		2851 => 32767,
		2852 => 32767,
		2853 => 32767,
		2854 => 32767,
		2855 => 32767,
		2856 => 32767,
		2857 => 32767,
		2858 => 32767,
		2859 => 32767,
		2860 => 32767,
		2861 => 32767,
		2862 => 32767,
		2863 => 32767,
		2864 => 32767,
		2865 => 32767,
		2866 => 32767,
		2867 => 32767,
		2868 => 32767,
		2869 => 32767,
		2870 => 32767,
		2871 => 32767,
		2872 => 32767,
		2873 => 32767,
		2874 => 32767,
		2875 => 32767,
		2876 => 32767,
		2877 => 32767,
		2878 => 32767,
		2879 => 32767,
		2880 => 32767,
		2881 => 32767,
		2882 => 32767,
		2883 => 32767,
		2884 => 32767,
		2885 => 32767,
		2886 => 32767,
		2887 => 32767,
		2888 => 32767,
		2889 => 32767,
		2890 => 32767,
		2891 => 32767,
		2892 => 32767,
		2893 => 32767,
		2894 => 32767,
		2895 => 32767,
		2896 => 32767,
		2897 => 32767,
		2898 => 32767,
		2899 => 32767,
		2900 => 32767,
		2901 => 32767,
		2902 => 32767,
		2903 => 32767,
		2904 => 32767,
		2905 => 32767,
		2906 => 32767,
		2907 => 32767,
		2908 => 32767,
		2909 => 32767,
		2910 => 32767,
		2911 => 32767,
		2912 => 32767,
		2913 => 32767,
		2914 => 32767,
		2915 => 32767,
		2916 => 32767,
		2917 => 32767,
		2918 => 32767,
		2919 => 32767,
		2920 => 32767,
		2921 => 32767,
		2922 => 32767,
		2923 => 32767,
		2924 => 32767,
		2925 => 32767,
		2926 => 32767,
		2927 => 32767,
		2928 => 32767,
		2929 => 32767,
		2930 => 32767,
		2931 => 32767,
		2932 => 32767,
		2933 => 32767,
		2934 => 32767,
		2935 => 32767,
		2936 => 32767,
		2937 => 32767,
		2938 => 32767,
		2939 => 32767,
		2940 => 32767,
		2941 => 32767,
		2942 => 32767,
		2943 => 32767,
		2944 => 32767,
		2945 => 32767,
		2946 => 32767,
		2947 => 32767,
		2948 => 32767,
		2949 => 32767,
		2950 => 32767,
		2951 => 32767,
		2952 => 32767,
		2953 => 32767,
		2954 => 32767,
		2955 => 32767,
		2956 => 32767,
		2957 => 32767,
		2958 => 32767,
		2959 => 32767,
		2960 => 32767,
		2961 => 32767,
		2962 => 32767,
		2963 => 32767,
		2964 => 32767,
		2965 => 32767,
		2966 => 32767,
		2967 => 32767,
		2968 => 32767,
		2969 => 32767,
		2970 => 32767,
		2971 => 32767,
		2972 => 32767,
		2973 => 32767,
		2974 => 32767,
		2975 => 32767,
		2976 => 32767,
		2977 => 32767,
		2978 => 32767,
		2979 => 32767,
		2980 => 32767,
		2981 => 32767,
		2982 => 32767,
		2983 => 32767,
		2984 => 32767,
		2985 => 32767,
		2986 => 32767,
		2987 => 32767,
		2988 => 32767,
		2989 => 32767,
		2990 => 32767,
		2991 => 32767,
		2992 => 32767,
		2993 => 32767,
		2994 => 32767,
		2995 => 32767,
		2996 => 32767,
		2997 => 32767,
		2998 => 32767,
		2999 => 32767,
		3000 => 32767,
		3001 => 32767,
		3002 => 32767,
		3003 => 32767,
		3004 => 32767,
		3005 => 32767,
		3006 => 32767,
		3007 => 32767,
		3008 => 32767,
		3009 => 32767,
		3010 => 32767,
		3011 => 32767,
		3012 => 32767,
		3013 => 32767,
		3014 => 32767,
		3015 => 32767,
		3016 => 32767,
		3017 => 32767,
		3018 => 32767,
		3019 => 32767,
		3020 => 32767,
		3021 => 32767,
		3022 => 32767,
		3023 => 32767,
		3024 => 32767,
		3025 => 32767,
		3026 => 32767,
		3027 => 32767,
		3028 => 32767,
		3029 => 32767,
		3030 => 32767,
		3031 => 32767,
		3032 => 32767,
		3033 => 32767,
		3034 => 32767,
		3035 => 32767,
		3036 => 32767,
		3037 => 32767,
		3038 => 32767,
		3039 => 32767,
		3040 => 32767,
		3041 => 32767,
		3042 => 32767,
		3043 => 32767,
		3044 => 32767,
		3045 => 32767,
		3046 => 32767,
		3047 => 32767,
		3048 => 32767,
		3049 => 32767,
		3050 => 32767,
		3051 => 32767,
		3052 => 32767,
		3053 => 32767,
		3054 => 32767,
		3055 => 32767,
		3056 => 32767,
		3057 => 32767,
		3058 => 32767,
		3059 => 32767,
		3060 => 32767,
		3061 => 32767,
		3062 => 32767,
		3063 => 32767,
		3064 => 32767,
		3065 => 32767,
		3066 => 32767,
		3067 => 32767,
		3068 => 32767,
		3069 => 32767,
		3070 => 32767,
		3071 => 32767,
		3072 => 32767,
		3073 => 32767,
		3074 => 32767,
		3075 => 32767,
		3076 => 32767,
		3077 => 32767,
		3078 => 32767,
		3079 => 32767,
		3080 => 32767,
		3081 => 32767,
		3082 => 32767,
		3083 => 32767,
		3084 => 32767,
		3085 => 32767,
		3086 => 32767,
		3087 => 32767,
		3088 => 32767,
		3089 => 32767,
		3090 => 32767,
		3091 => 32767,
		3092 => 32767,
		3093 => 32767,
		3094 => 32767,
		3095 => 32767,
		3096 => 32767,
		3097 => 32767,
		3098 => 32767,
		3099 => 32767,
		3100 => 32767,
		3101 => 32767,
		3102 => 32767,
		3103 => 32767,
		3104 => 32767,
		3105 => 32767,
		3106 => 32767,
		3107 => 32767,
		3108 => 32767,
		3109 => 32767,
		3110 => 32767,
		3111 => 32767,
		3112 => 32767,
		3113 => 32767,
		3114 => 32767,
		3115 => 32767,
		3116 => 32767,
		3117 => 32767,
		3118 => 32767,
		3119 => 32767,
		3120 => 32767,
		3121 => 32767,
		3122 => 32767,
		3123 => 32767,
		3124 => 32767,
		3125 => 32767,
		3126 => 32767,
		3127 => 32767,
		3128 => 32767,
		3129 => 32767,
		3130 => 32767,
		3131 => 32767,
		3132 => 32767,
		3133 => 32767,
		3134 => 32767,
		3135 => 32767,
		3136 => 32767,
		3137 => 32767,
		3138 => 32767,
		3139 => 32767,
		3140 => 32767,
		3141 => 32767,
		3142 => 32767,
		3143 => 32767,
		3144 => 32767,
		3145 => 32767,
		3146 => 32767,
		3147 => 32767,
		3148 => 32767,
		3149 => 32767,
		3150 => 32767,
		3151 => 32767,
		3152 => 32767,
		3153 => 32767,
		3154 => 32767,
		3155 => 32767,
		3156 => 32767,
		3157 => 32767,
		3158 => 32767,
		3159 => 32767,
		3160 => 32767,
		3161 => 32767,
		3162 => 32767,
		3163 => 32767,
		3164 => 32767,
		3165 => 32767,
		3166 => 32767,
		3167 => 32767,
		3168 => 32767,
		3169 => 32767,
		3170 => 32767,
		3171 => 32767,
		3172 => 32767,
		3173 => 32767,
		3174 => 32767,
		3175 => 32767,
		3176 => 32767,
		3177 => 32767,
		3178 => 32767,
		3179 => 32767,
		3180 => 32767,
		3181 => 32767,
		3182 => 32767,
		3183 => 32767,
		3184 => 32767,
		3185 => 32767,
		3186 => 32767,
		3187 => 32767,
		3188 => 32767,
		3189 => 32767,
		3190 => 32767,
		3191 => 32767,
		3192 => 32767,
		3193 => 32767,
		3194 => 32767,
		3195 => 32767,
		3196 => 32767,
		3197 => 32767,
		3198 => 32767,
		3199 => 32767,
		3200 => 32767,
		3201 => 32767,
		3202 => 32767,
		3203 => 32767,
		3204 => 32767,
		3205 => 32767,
		3206 => 32767,
		3207 => 32767,
		3208 => 32767,
		3209 => 32767,
		3210 => 32767,
		3211 => 32767,
		3212 => 32767,
		3213 => 32767,
		3214 => 32767,
		3215 => 32767,
		3216 => 32767,
		3217 => 32767,
		3218 => 32767,
		3219 => 32767,
		3220 => 32767,
		3221 => 32767,
		3222 => 32767,
		3223 => 32767,
		3224 => 32767,
		3225 => 32767,
		3226 => 32767,
		3227 => 32767,
		3228 => 32767,
		3229 => 32767,
		3230 => 32767,
		3231 => 32767,
		3232 => 32767,
		3233 => 32767,
		3234 => 32767,
		3235 => 32767,
		3236 => 32767,
		3237 => 32767,
		3238 => 32767,
		3239 => 32767,
		3240 => 32767,
		3241 => 32767,
		3242 => 32767,
		3243 => 32767,
		3244 => 32767,
		3245 => 32767,
		3246 => 32767,
		3247 => 32767,
		3248 => 32767,
		3249 => 32767,
		3250 => 32767,
		3251 => 32767,
		3252 => 32767,
		3253 => 32767,
		3254 => 32767,
		3255 => 32767,
		3256 => 32767,
		3257 => 32767,
		3258 => 32767,
		3259 => 32767,
		3260 => 32767,
		3261 => 32767,
		3262 => 32767,
		3263 => 32767,
		3264 => 32767,
		3265 => 32767,
		3266 => 32767,
		3267 => 32767,
		3268 => 32767,
		3269 => 32767,
		3270 => 32767,
		3271 => 32767,
		3272 => 32767,
		3273 => 32767,
		3274 => 32767,
		3275 => 32767,
		3276 => 32767,
		3277 => 32767,
		3278 => 32767,
		3279 => 32767,
		3280 => 32767,
		3281 => 32767,
		3282 => 32767,
		3283 => 32767,
		3284 => 32767,
		3285 => 32767,
		3286 => 32767,
		3287 => 32767,
		3288 => 32767,
		3289 => 32767,
		3290 => 32767,
		3291 => 32767,
		3292 => 32767,
		3293 => 32767,
		3294 => 32767,
		3295 => 32767,
		3296 => 32767,
		3297 => 32767,
		3298 => 32767,
		3299 => 32767,
		3300 => 32767,
		3301 => 32767,
		3302 => 32767,
		3303 => 32767,
		3304 => 32767,
		3305 => 32767,
		3306 => 32767,
		3307 => 32767,
		3308 => 32767,
		3309 => 32767,
		3310 => 32767,
		3311 => 32767,
		3312 => 32767,
		3313 => 32767,
		3314 => 32767,
		3315 => 32767,
		3316 => 32767,
		3317 => 32767,
		3318 => 32767,
		3319 => 32767,
		3320 => 32767,
		3321 => 32767,
		3322 => 32767,
		3323 => 32767,
		3324 => 32767,
		3325 => 32767,
		3326 => 32767,
		3327 => 32767,
		3328 => 32767,
		3329 => 32767,
		3330 => 32767,
		3331 => 32767,
		3332 => 32767,
		3333 => 32767,
		3334 => 32767,
		3335 => 32767,
		3336 => 32767,
		3337 => 32767,
		3338 => 32767,
		3339 => 32767,
		3340 => 32767,
		3341 => 32767,
		3342 => 32767,
		3343 => 32767,
		3344 => 32767,
		3345 => 32767,
		3346 => 32767,
		3347 => 32767,
		3348 => 32767,
		3349 => 32767,
		3350 => 32767,
		3351 => 32767,
		3352 => 32767,
		3353 => 32767,
		3354 => 32767,
		3355 => 32767,
		3356 => 32767,
		3357 => 32767,
		3358 => 32767,
		3359 => 32767,
		3360 => 32767,
		3361 => 32767,
		3362 => 32767,
		3363 => 32767,
		3364 => 32767,
		3365 => 32767,
		3366 => 32767,
		3367 => 32767,
		3368 => 32767,
		3369 => 32767,
		3370 => 32767,
		3371 => 32767,
		3372 => 32767,
		3373 => 32767,
		3374 => 32767,
		3375 => 32767,
		3376 => 32767,
		3377 => 32767,
		3378 => 32767,
		3379 => 32767,
		3380 => 32767,
		3381 => 32767,
		3382 => 32767,
		3383 => 32767,
		3384 => 32767,
		3385 => 32767,
		3386 => 32767,
		3387 => 32767,
		3388 => 32767,
		3389 => 32767,
		3390 => 32767,
		3391 => 32767,
		3392 => 32767,
		3393 => 32767,
		3394 => 32767,
		3395 => 32767,
		3396 => 32767,
		3397 => 32767,
		3398 => 32767,
		3399 => 32767,
		3400 => 32767,
		3401 => 32767,
		3402 => 32767,
		3403 => 32767,
		3404 => 32767,
		3405 => 32767,
		3406 => 32767,
		3407 => 32767,
		3408 => 32767,
		3409 => 32767,
		3410 => 32767,
		3411 => 32767,
		3412 => 32767,
		3413 => 32767,
		3414 => 32767,
		3415 => 32767,
		3416 => 32767,
		3417 => 32767,
		3418 => 32767,
		3419 => 32767,
		3420 => 32767,
		3421 => 32767,
		3422 => 32767,
		3423 => 32767,
		3424 => 32767,
		3425 => 32767,
		3426 => 32767,
		3427 => 32767,
		3428 => 32767,
		3429 => 32767,
		3430 => 32767,
		3431 => 32767,
		3432 => 32767,
		3433 => 32767,
		3434 => 32767,
		3435 => 32767,
		3436 => 32767,
		3437 => 32767,
		3438 => 32767,
		3439 => 32767,
		3440 => 32767,
		3441 => 32767,
		3442 => 32767,
		3443 => 32767,
		3444 => 32767,
		3445 => 32767,
		3446 => 32767,
		3447 => 32767,
		3448 => 32767,
		3449 => 32767,
		3450 => 32767,
		3451 => 32767,
		3452 => 32767,
		3453 => 32767,
		3454 => 32767,
		3455 => 32767,
		3456 => 32767,
		3457 => 32767,
		3458 => 32767,
		3459 => 32767,
		3460 => 32767,
		3461 => 32767,
		3462 => 32767,
		3463 => 32767,
		3464 => 32767,
		3465 => 32767,
		3466 => 32767,
		3467 => 32767,
		3468 => 32767,
		3469 => 32767,
		3470 => 32767,
		3471 => 32767,
		3472 => 32767,
		3473 => 32767,
		3474 => 32767,
		3475 => 32767,
		3476 => 32767,
		3477 => 32767,
		3478 => 32767,
		3479 => 32767,
		3480 => 32767,
		3481 => 32767,
		3482 => 32767,
		3483 => 32767,
		3484 => 32767,
		3485 => 32767,
		3486 => 32767,
		3487 => 32767,
		3488 => 32767,
		3489 => 32767,
		3490 => 32767,
		3491 => 32767,
		3492 => 32767,
		3493 => 32767,
		3494 => 32767,
		3495 => 32767,
		3496 => 32767,
		3497 => 32767,
		3498 => 32767,
		3499 => 32767,
		3500 => 32767,
		3501 => 32767,
		3502 => 32767,
		3503 => 32767,
		3504 => 32767,
		3505 => 32767,
		3506 => 32767,
		3507 => 32767,
		3508 => 32767,
		3509 => 32767,
		3510 => 32767,
		3511 => 32767,
		3512 => 32767,
		3513 => 32767,
		3514 => 32767,
		3515 => 32767,
		3516 => 32767,
		3517 => 32767,
		3518 => 32767,
		3519 => 32767,
		3520 => 32767,
		3521 => 32767,
		3522 => 32767,
		3523 => 32767,
		3524 => 32767,
		3525 => 32767,
		3526 => 32767,
		3527 => 32767,
		3528 => 32767,
		3529 => 32767,
		3530 => 32767,
		3531 => 32767,
		3532 => 32767,
		3533 => 32767,
		3534 => 32767,
		3535 => 32767,
		3536 => 32767,
		3537 => 32767,
		3538 => 32767,
		3539 => 32767,
		3540 => 32767,
		3541 => 32767,
		3542 => 32767,
		3543 => 32767,
		3544 => 32767,
		3545 => 32767,
		3546 => 32767,
		3547 => 32767,
		3548 => 32767,
		3549 => 32767,
		3550 => 32767,
		3551 => 32767,
		3552 => 32767,
		3553 => 32767,
		3554 => 32767,
		3555 => 32767,
		3556 => 32767,
		3557 => 32767,
		3558 => 32767,
		3559 => 32767,
		3560 => 32767,
		3561 => 32767,
		3562 => 32767,
		3563 => 32767,
		3564 => 32767,
		3565 => 32767,
		3566 => 32767,
		3567 => 32767,
		3568 => 32767,
		3569 => 32767,
		3570 => 32767,
		3571 => 32767,
		3572 => 32767,
		3573 => 32767,
		3574 => 32767,
		3575 => 32767,
		3576 => 32767,
		3577 => 32767,
		3578 => 32767,
		3579 => 32767,
		3580 => 32767,
		3581 => 32767,
		3582 => 32767,
		3583 => 32767,
		3584 => 32767,
		3585 => 32767,
		3586 => 32767,
		3587 => 32767,
		3588 => 32767,
		3589 => 32767,
		3590 => 32767,
		3591 => 32767,
		3592 => 32767,
		3593 => 32767,
		3594 => 32767,
		3595 => 32767,
		3596 => 32767,
		3597 => 32767,
		3598 => 32767,
		3599 => 32767,
		3600 => 32767,
		3601 => 32767,
		3602 => 32767,
		3603 => 32767,
		3604 => 32767,
		3605 => 32767,
		3606 => 32767,
		3607 => 32767,
		3608 => 32767,
		3609 => 32767,
		3610 => 32767,
		3611 => 32767,
		3612 => 32767,
		3613 => 32767,
		3614 => 32767,
		3615 => 32767,
		3616 => 32767,
		3617 => 32767,
		3618 => 32767,
		3619 => 32767,
		3620 => 32767,
		3621 => 32767,
		3622 => 32767,
		3623 => 32767,
		3624 => 32767,
		3625 => 32767,
		3626 => 32767,
		3627 => 32767,
		3628 => 32767,
		3629 => 32767,
		3630 => 32767,
		3631 => 32767,
		3632 => 32767,
		3633 => 32767,
		3634 => 32767,
		3635 => 32767,
		3636 => 32767,
		3637 => 32767,
		3638 => 32767,
		3639 => 32767,
		3640 => 32767,
		3641 => 32767,
		3642 => 32767,
		3643 => 32767,
		3644 => 32767,
		3645 => 32767,
		3646 => 32767,
		3647 => 32767,
		3648 => 32767,
		3649 => 32767,
		3650 => 32767,
		3651 => 32767,
		3652 => 32767,
		3653 => 32767,
		3654 => 32767,
		3655 => 32767,
		3656 => 32767,
		3657 => 32767,
		3658 => 32767,
		3659 => 32767,
		3660 => 32767,
		3661 => 32767,
		3662 => 32767,
		3663 => 32767,
		3664 => 32767,
		3665 => 32767,
		3666 => 32767,
		3667 => 32767,
		3668 => 32767,
		3669 => 32767,
		3670 => 32767,
		3671 => 32767,
		3672 => 32767,
		3673 => 32767,
		3674 => 32767,
		3675 => 32767,
		3676 => 32767,
		3677 => 32767,
		3678 => 32767,
		3679 => 32767,
		3680 => 32767,
		3681 => 32767,
		3682 => 32767,
		3683 => 32767,
		3684 => 32767,
		3685 => 32767,
		3686 => 32767,
		3687 => 32767,
		3688 => 32767,
		3689 => 32767,
		3690 => 32767,
		3691 => 32767,
		3692 => 32767,
		3693 => 32767,
		3694 => 32767,
		3695 => 32767,
		3696 => 32767,
		3697 => 32767,
		3698 => 32767,
		3699 => 32767,
		3700 => 32767,
		3701 => 32767,
		3702 => 32767,
		3703 => 32767,
		3704 => 32767,
		3705 => 32767,
		3706 => 32767,
		3707 => 32767,
		3708 => 32767,
		3709 => 32767,
		3710 => 32767,
		3711 => 32767,
		3712 => 32767,
		3713 => 32767,
		3714 => 32767,
		3715 => 32767,
		3716 => 32767,
		3717 => 32767,
		3718 => 32767,
		3719 => 32767,
		3720 => 32767,
		3721 => 32767,
		3722 => 32767,
		3723 => 32767,
		3724 => 32767,
		3725 => 32767,
		3726 => 32767,
		3727 => 32767,
		3728 => 32767,
		3729 => 32767,
		3730 => 32767,
		3731 => 32767,
		3732 => 32767,
		3733 => 32767,
		3734 => 32767,
		3735 => 32767,
		3736 => 32767,
		3737 => 32767,
		3738 => 32767,
		3739 => 32767,
		3740 => 32767,
		3741 => 32767,
		3742 => 32767,
		3743 => 32767,
		3744 => 32767,
		3745 => 32767,
		3746 => 32767,
		3747 => 32767,
		3748 => 32767,
		3749 => 32767,
		3750 => 32767,
		3751 => 32767,
		3752 => 32767,
		3753 => 32767,
		3754 => 32767,
		3755 => 32767,
		3756 => 32767,
		3757 => 32767,
		3758 => 32767,
		3759 => 32767,
		3760 => 32767,
		3761 => 32767,
		3762 => 32767,
		3763 => 32767,
		3764 => 32767,
		3765 => 32767,
		3766 => 32767,
		3767 => 32767,
		3768 => 32767,
		3769 => 32767,
		3770 => 32767,
		3771 => 32767,
		3772 => 32767,
		3773 => 32767,
		3774 => 32767,
		3775 => 32767,
		3776 => 32767,
		3777 => 32767,
		3778 => 32767,
		3779 => 32767,
		3780 => 32767,
		3781 => 32767,
		3782 => 32767,
		3783 => 32767,
		3784 => 32767,
		3785 => 32767,
		3786 => 32767,
		3787 => 32767,
		3788 => 32767,
		3789 => 32767,
		3790 => 32767,
		3791 => 32767,
		3792 => 32767,
		3793 => 32767,
		3794 => 32767,
		3795 => 32767,
		3796 => 32767,
		3797 => 32767,
		3798 => 32767,
		3799 => 32767,
		3800 => 32767,
		3801 => 32767,
		3802 => 32767,
		3803 => 32767,
		3804 => 32767,
		3805 => 32767,
		3806 => 32767,
		3807 => 32767,
		3808 => 32767,
		3809 => 32767,
		3810 => 32767,
		3811 => 32767,
		3812 => 32767,
		3813 => 32767,
		3814 => 32767,
		3815 => 32767,
		3816 => 32767,
		3817 => 32767,
		3818 => 32767,
		3819 => 32767,
		3820 => 32767,
		3821 => 32767,
		3822 => 32767,
		3823 => 32767,
		3824 => 32767,
		3825 => 32767,
		3826 => 32767,
		3827 => 32767,
		3828 => 32767,
		3829 => 32767,
		3830 => 32767,
		3831 => 32767,
		3832 => 32767,
		3833 => 32767,
		3834 => 32767,
		3835 => 32767,
		3836 => 32767,
		3837 => 32767,
		3838 => 32767,
		3839 => 32767,
		3840 => 32767,
		3841 => 32767,
		3842 => 32767,
		3843 => 32767,
		3844 => 32767,
		3845 => 32767,
		3846 => 32767,
		3847 => 32767,
		3848 => 32767,
		3849 => 32767,
		3850 => 32767,
		3851 => 32767,
		3852 => 32767,
		3853 => 32767,
		3854 => 32767,
		3855 => 32767,
		3856 => 32767,
		3857 => 32767,
		3858 => 32767,
		3859 => 32767,
		3860 => 32767,
		3861 => 32767,
		3862 => 32767,
		3863 => 32767,
		3864 => 32767,
		3865 => 32767,
		3866 => 32767,
		3867 => 32767,
		3868 => 32767,
		3869 => 32767,
		3870 => 32767,
		3871 => 32767,
		3872 => 32767,
		3873 => 32767,
		3874 => 32767,
		3875 => 32767,
		3876 => 32767,
		3877 => 32767,
		3878 => 32767,
		3879 => 32767,
		3880 => 32767,
		3881 => 32767,
		3882 => 32767,
		3883 => 32767,
		3884 => 32767,
		3885 => 32767,
		3886 => 32767,
		3887 => 32767,
		3888 => 32767,
		3889 => 32767,
		3890 => 32767,
		3891 => 32767,
		3892 => 32767,
		3893 => 32767,
		3894 => 32767,
		3895 => 32767,
		3896 => 32767,
		3897 => 32767,
		3898 => 32767,
		3899 => 32767,
		3900 => 32767,
		3901 => 32767,
		3902 => 32767,
		3903 => 32767,
		3904 => 32767,
		3905 => 32767,
		3906 => 32767,
		3907 => 32767,
		3908 => 32767,
		3909 => 32767,
		3910 => 32767,
		3911 => 32767,
		3912 => 32767,
		3913 => 32767,
		3914 => 32767,
		3915 => 32767,
		3916 => 32767,
		3917 => 32767,
		3918 => 32767,
		3919 => 32767,
		3920 => 32767,
		3921 => 32767,
		3922 => 32767,
		3923 => 32767,
		3924 => 32767,
		3925 => 32767,
		3926 => 32767,
		3927 => 32767,
		3928 => 32767,
		3929 => 32767,
		3930 => 32767,
		3931 => 32767,
		3932 => 32767,
		3933 => 32767,
		3934 => 32767,
		3935 => 32767,
		3936 => 32767,
		3937 => 32767,
		3938 => 32767,
		3939 => 32767,
		3940 => 32767,
		3941 => 32767,
		3942 => 32767,
		3943 => 32767,
		3944 => 32767,
		3945 => 32767,
		3946 => 32767,
		3947 => 32767,
		3948 => 32767,
		3949 => 32767,
		3950 => 32767,
		3951 => 32767,
		3952 => 32767,
		3953 => 32767,
		3954 => 32767,
		3955 => 32767,
		3956 => 32767,
		3957 => 32767,
		3958 => 32767,
		3959 => 32767,
		3960 => 32767,
		3961 => 32767,
		3962 => 32767,
		3963 => 32767,
		3964 => 32767,
		3965 => 32767,
		3966 => 32767,
		3967 => 32767,
		3968 => 32767,
		3969 => 32767,
		3970 => 32767,
		3971 => 32767,
		3972 => 32767,
		3973 => 32767,
		3974 => 32767,
		3975 => 32767,
		3976 => 32767,
		3977 => 32767,
		3978 => 32767,
		3979 => 32767,
		3980 => 32767,
		3981 => 32767,
		3982 => 32767,
		3983 => 32767,
		3984 => 32767,
		3985 => 32767,
		3986 => 32767,
		3987 => 32767,
		3988 => 32767,
		3989 => 32767,
		3990 => 32767,
		3991 => 32767,
		3992 => 32767,
		3993 => 32767,
		3994 => 32767,
		3995 => 32767,
		3996 => 32767,
		3997 => 32767,
		3998 => 32767,
		3999 => 32767,
		4000 => 32767,
		4001 => 32767,
		4002 => 32767,
		4003 => 32767,
		4004 => 32767,
		4005 => 32767,
		4006 => 32767,
		4007 => 32767,
		4008 => 32767,
		4009 => 32767,
		4010 => 32767,
		4011 => 32767,
		4012 => 32767,
		4013 => 32767,
		4014 => 32767,
		4015 => 32767,
		4016 => 32767,
		4017 => 32767,
		4018 => 32767,
		4019 => 32767,
		4020 => 32767,
		4021 => 32767,
		4022 => 32767,
		4023 => 32767,
		4024 => 32767,
		4025 => 32767,
		4026 => 32767,
		4027 => 32767,
		4028 => 32767,
		4029 => 32767,
		4030 => 32767,
		4031 => 32767,
		4032 => 32767,
		4033 => 32767,
		4034 => 32767,
		4035 => 32767,
		4036 => 32767,
		4037 => 32767,
		4038 => 32767,
		4039 => 32767,
		4040 => 32767,
		4041 => 32767,
		4042 => 32767,
		4043 => 32767,
		4044 => 32767,
		4045 => 32767,
		4046 => 32767,
		4047 => 32767,
		4048 => 32767,
		4049 => 32767,
		4050 => 32767,
		4051 => 32767,
		4052 => 32767,
		4053 => 32767,
		4054 => 32767,
		4055 => 32767,
		4056 => 32767,
		4057 => 32767,
		4058 => 32767,
		4059 => 32767,
		4060 => 32767,
		4061 => 32767,
		4062 => 32767,
		4063 => 32767,
		4064 => 32767,
		4065 => 32767,
		4066 => 32767,
		4067 => 32767,
		4068 => 32767,
		4069 => 32767,
		4070 => 32767,
		4071 => 32767,
		4072 => 32767,
		4073 => 32767,
		4074 => 32767,
		4075 => 32767,
		4076 => 32767,
		4077 => 32767,
		4078 => 32767,
		4079 => 32767,
		4080 => 32767,
		4081 => 32767,
		4082 => 32767,
		4083 => 32767,
		4084 => 32767,
		4085 => 32767,
		4086 => 32767,
		4087 => 32767,
		4088 => 32767,
		4089 => 32767,
		4090 => 32767,
		4091 => 32767,
		4092 => 32767,
		4093 => 32767,
		4094 => 32767,
		4095 => 32767
);

begin
	sigmoid_out <= std_logic_vector(TO_SIGNED(LUT(TO_INTEGER(unsigned(address))),16));
end beh;
