library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LUT_4096 is
	port (
		address : in  std_logic_vector(12 downto 0);
		dds_out : out std_logic_vector(15 downto 0) 
	);
end LUT_4096;

architecture beh of LUT_4096 is
	type LUT_t is array (natural range 0 to 4095) of integer;
	constant LUT: LUT_t := (
		0 => 16384,
		1 => 16406,
		2 => 16428,
		3 => 16450,
		4 => 16472,
		5 => 16494,
		6 => 16516,
		7 => 16538,
		8 => 16560,
		9 => 16582,
		10 => 16604,
		11 => 16626,
		12 => 16648,
		13 => 16670,
		14 => 16692,
		15 => 16714,
		16 => 16736,
		17 => 16758,
		18 => 16780,
		19 => 16801,
		20 => 16823,
		21 => 16845,
		22 => 16867,
		23 => 16889,
		24 => 16911,
		25 => 16933,
		26 => 16955,
		27 => 16977,
		28 => 16999,
		29 => 17021,
		30 => 17043,
		31 => 17065,
		32 => 17087,
		33 => 17109,
		34 => 17131,
		35 => 17153,
		36 => 17175,
		37 => 17197,
		38 => 17219,
		39 => 17241,
		40 => 17263,
		41 => 17285,
		42 => 17307,
		43 => 17329,
		44 => 17351,
		45 => 17373,
		46 => 17394,
		47 => 17416,
		48 => 17438,
		49 => 17460,
		50 => 17482,
		51 => 17504,
		52 => 17526,
		53 => 17548,
		54 => 17570,
		55 => 17592,
		56 => 17613,
		57 => 17635,
		58 => 17657,
		59 => 17679,
		60 => 17701,
		61 => 17723,
		62 => 17745,
		63 => 17766,
		64 => 17788,
		65 => 17810,
		66 => 17832,
		67 => 17854,
		68 => 17876,
		69 => 17897,
		70 => 17919,
		71 => 17941,
		72 => 17963,
		73 => 17985,
		74 => 18007,
		75 => 18028,
		76 => 18050,
		77 => 18072,
		78 => 18094,
		79 => 18115,
		80 => 18137,
		81 => 18159,
		82 => 18181,
		83 => 18202,
		84 => 18224,
		85 => 18246,
		86 => 18268,
		87 => 18289,
		88 => 18311,
		89 => 18333,
		90 => 18354,
		91 => 18376,
		92 => 18398,
		93 => 18419,
		94 => 18441,
		95 => 18463,
		96 => 18484,
		97 => 18506,
		98 => 18528,
		99 => 18549,
		100 => 18571,
		101 => 18592,
		102 => 18614,
		103 => 18636,
		104 => 18657,
		105 => 18679,
		106 => 18700,
		107 => 18722,
		108 => 18743,
		109 => 18765,
		110 => 18787,
		111 => 18808,
		112 => 18830,
		113 => 18851,
		114 => 18873,
		115 => 18894,
		116 => 18916,
		117 => 18937,
		118 => 18959,
		119 => 18980,
		120 => 19001,
		121 => 19023,
		122 => 19044,
		123 => 19066,
		124 => 19087,
		125 => 19109,
		126 => 19130,
		127 => 19151,
		128 => 19173,
		129 => 19194,
		130 => 19215,
		131 => 19237,
		132 => 19258,
		133 => 19279,
		134 => 19301,
		135 => 19322,
		136 => 19343,
		137 => 19365,
		138 => 19386,
		139 => 19407,
		140 => 19428,
		141 => 19450,
		142 => 19471,
		143 => 19492,
		144 => 19513,
		145 => 19534,
		146 => 19556,
		147 => 19577,
		148 => 19598,
		149 => 19619,
		150 => 19640,
		151 => 19661,
		152 => 19683,
		153 => 19704,
		154 => 19725,
		155 => 19746,
		156 => 19767,
		157 => 19788,
		158 => 19809,
		159 => 19830,
		160 => 19851,
		161 => 19872,
		162 => 19893,
		163 => 19914,
		164 => 19935,
		165 => 19956,
		166 => 19977,
		167 => 19998,
		168 => 20019,
		169 => 20040,
		170 => 20061,
		171 => 20082,
		172 => 20102,
		173 => 20123,
		174 => 20144,
		175 => 20165,
		176 => 20186,
		177 => 20207,
		178 => 20227,
		179 => 20248,
		180 => 20269,
		181 => 20290,
		182 => 20310,
		183 => 20331,
		184 => 20352,
		185 => 20373,
		186 => 20393,
		187 => 20414,
		188 => 20435,
		189 => 20455,
		190 => 20476,
		191 => 20497,
		192 => 20517,
		193 => 20538,
		194 => 20558,
		195 => 20579,
		196 => 20599,
		197 => 20620,
		198 => 20641,
		199 => 20661,
		200 => 20682,
		201 => 20702,
		202 => 20723,
		203 => 20743,
		204 => 20763,
		205 => 20784,
		206 => 20804,
		207 => 20825,
		208 => 20845,
		209 => 20865,
		210 => 20886,
		211 => 20906,
		212 => 20926,
		213 => 20947,
		214 => 20967,
		215 => 20987,
		216 => 21008,
		217 => 21028,
		218 => 21048,
		219 => 21068,
		220 => 21088,
		221 => 21109,
		222 => 21129,
		223 => 21149,
		224 => 21169,
		225 => 21189,
		226 => 21209,
		227 => 21229,
		228 => 21249,
		229 => 21269,
		230 => 21290,
		231 => 21310,
		232 => 21330,
		233 => 21350,
		234 => 21370,
		235 => 21389,
		236 => 21409,
		237 => 21429,
		238 => 21449,
		239 => 21469,
		240 => 21489,
		241 => 21509,
		242 => 21529,
		243 => 21549,
		244 => 21568,
		245 => 21588,
		246 => 21608,
		247 => 21628,
		248 => 21647,
		249 => 21667,
		250 => 21687,
		251 => 21707,
		252 => 21726,
		253 => 21746,
		254 => 21766,
		255 => 21785,
		256 => 21805,
		257 => 21824,
		258 => 21844,
		259 => 21863,
		260 => 21883,
		261 => 21902,
		262 => 21922,
		263 => 21941,
		264 => 21961,
		265 => 21980,
		266 => 22000,
		267 => 22019,
		268 => 22039,
		269 => 22058,
		270 => 22077,
		271 => 22097,
		272 => 22116,
		273 => 22135,
		274 => 22155,
		275 => 22174,
		276 => 22193,
		277 => 22212,
		278 => 22232,
		279 => 22251,
		280 => 22270,
		281 => 22289,
		282 => 22308,
		283 => 22327,
		284 => 22346,
		285 => 22365,
		286 => 22385,
		287 => 22404,
		288 => 22423,
		289 => 22442,
		290 => 22461,
		291 => 22480,
		292 => 22499,
		293 => 22517,
		294 => 22536,
		295 => 22555,
		296 => 22574,
		297 => 22593,
		298 => 22612,
		299 => 22631,
		300 => 22649,
		301 => 22668,
		302 => 22687,
		303 => 22706,
		304 => 22724,
		305 => 22743,
		306 => 22762,
		307 => 22780,
		308 => 22799,
		309 => 22818,
		310 => 22836,
		311 => 22855,
		312 => 22873,
		313 => 22892,
		314 => 22911,
		315 => 22929,
		316 => 22948,
		317 => 22966,
		318 => 22984,
		319 => 23003,
		320 => 23021,
		321 => 23040,
		322 => 23058,
		323 => 23076,
		324 => 23095,
		325 => 23113,
		326 => 23131,
		327 => 23149,
		328 => 23168,
		329 => 23186,
		330 => 23204,
		331 => 23222,
		332 => 23241,
		333 => 23259,
		334 => 23277,
		335 => 23295,
		336 => 23313,
		337 => 23331,
		338 => 23349,
		339 => 23367,
		340 => 23385,
		341 => 23403,
		342 => 23421,
		343 => 23439,
		344 => 23457,
		345 => 23475,
		346 => 23493,
		347 => 23510,
		348 => 23528,
		349 => 23546,
		350 => 23564,
		351 => 23582,
		352 => 23599,
		353 => 23617,
		354 => 23635,
		355 => 23652,
		356 => 23670,
		357 => 23688,
		358 => 23705,
		359 => 23723,
		360 => 23741,
		361 => 23758,
		362 => 23776,
		363 => 23793,
		364 => 23811,
		365 => 23828,
		366 => 23846,
		367 => 23863,
		368 => 23880,
		369 => 23898,
		370 => 23915,
		371 => 23933,
		372 => 23950,
		373 => 23967,
		374 => 23984,
		375 => 24002,
		376 => 24019,
		377 => 24036,
		378 => 24053,
		379 => 24071,
		380 => 24088,
		381 => 24105,
		382 => 24122,
		383 => 24139,
		384 => 24156,
		385 => 24173,
		386 => 24190,
		387 => 24207,
		388 => 24224,
		389 => 24241,
		390 => 24258,
		391 => 24275,
		392 => 24292,
		393 => 24309,
		394 => 24325,
		395 => 24342,
		396 => 24359,
		397 => 24376,
		398 => 24393,
		399 => 24409,
		400 => 24426,
		401 => 24443,
		402 => 24459,
		403 => 24476,
		404 => 24493,
		405 => 24509,
		406 => 24526,
		407 => 24542,
		408 => 24559,
		409 => 24576,
		410 => 24592,
		411 => 24608,
		412 => 24625,
		413 => 24641,
		414 => 24658,
		415 => 24674,
		416 => 24691,
		417 => 24707,
		418 => 24723,
		419 => 24739,
		420 => 24756,
		421 => 24772,
		422 => 24788,
		423 => 24804,
		424 => 24821,
		425 => 24837,
		426 => 24853,
		427 => 24869,
		428 => 24885,
		429 => 24901,
		430 => 24917,
		431 => 24933,
		432 => 24949,
		433 => 24965,
		434 => 24981,
		435 => 24997,
		436 => 25013,
		437 => 25029,
		438 => 25045,
		439 => 25061,
		440 => 25076,
		441 => 25092,
		442 => 25108,
		443 => 25124,
		444 => 25139,
		445 => 25155,
		446 => 25171,
		447 => 25187,
		448 => 25202,
		449 => 25218,
		450 => 25233,
		451 => 25249,
		452 => 25264,
		453 => 25280,
		454 => 25296,
		455 => 25311,
		456 => 25326,
		457 => 25342,
		458 => 25357,
		459 => 25373,
		460 => 25388,
		461 => 25403,
		462 => 25419,
		463 => 25434,
		464 => 25449,
		465 => 25465,
		466 => 25480,
		467 => 25495,
		468 => 25510,
		469 => 25525,
		470 => 25541,
		471 => 25556,
		472 => 25571,
		473 => 25586,
		474 => 25601,
		475 => 25616,
		476 => 25631,
		477 => 25646,
		478 => 25661,
		479 => 25676,
		480 => 25691,
		481 => 25706,
		482 => 25720,
		483 => 25735,
		484 => 25750,
		485 => 25765,
		486 => 25780,
		487 => 25794,
		488 => 25809,
		489 => 25824,
		490 => 25839,
		491 => 25853,
		492 => 25868,
		493 => 25883,
		494 => 25897,
		495 => 25912,
		496 => 25926,
		497 => 25941,
		498 => 25955,
		499 => 25970,
		500 => 25984,
		501 => 25999,
		502 => 26013,
		503 => 26027,
		504 => 26042,
		505 => 26056,
		506 => 26070,
		507 => 26085,
		508 => 26099,
		509 => 26113,
		510 => 26128,
		511 => 26142,
		512 => 26156,
		513 => 26170,
		514 => 26184,
		515 => 26198,
		516 => 26212,
		517 => 26227,
		518 => 26241,
		519 => 26255,
		520 => 26269,
		521 => 26283,
		522 => 26297,
		523 => 26311,
		524 => 26324,
		525 => 26338,
		526 => 26352,
		527 => 26366,
		528 => 26380,
		529 => 26394,
		530 => 26407,
		531 => 26421,
		532 => 26435,
		533 => 26449,
		534 => 26462,
		535 => 26476,
		536 => 26490,
		537 => 26503,
		538 => 26517,
		539 => 26530,
		540 => 26544,
		541 => 26558,
		542 => 26571,
		543 => 26585,
		544 => 26598,
		545 => 26611,
		546 => 26625,
		547 => 26638,
		548 => 26652,
		549 => 26665,
		550 => 26678,
		551 => 26692,
		552 => 26705,
		553 => 26718,
		554 => 26731,
		555 => 26745,
		556 => 26758,
		557 => 26771,
		558 => 26784,
		559 => 26797,
		560 => 26810,
		561 => 26823,
		562 => 26836,
		563 => 26849,
		564 => 26863,
		565 => 26876,
		566 => 26888,
		567 => 26901,
		568 => 26914,
		569 => 26927,
		570 => 26940,
		571 => 26953,
		572 => 26966,
		573 => 26979,
		574 => 26991,
		575 => 27004,
		576 => 27017,
		577 => 27030,
		578 => 27042,
		579 => 27055,
		580 => 27068,
		581 => 27080,
		582 => 27093,
		583 => 27106,
		584 => 27118,
		585 => 27131,
		586 => 27143,
		587 => 27156,
		588 => 27168,
		589 => 27181,
		590 => 27193,
		591 => 27205,
		592 => 27218,
		593 => 27230,
		594 => 27243,
		595 => 27255,
		596 => 27267,
		597 => 27280,
		598 => 27292,
		599 => 27304,
		600 => 27316,
		601 => 27328,
		602 => 27341,
		603 => 27353,
		604 => 27365,
		605 => 27377,
		606 => 27389,
		607 => 27401,
		608 => 27413,
		609 => 27425,
		610 => 27437,
		611 => 27449,
		612 => 27461,
		613 => 27473,
		614 => 27485,
		615 => 27497,
		616 => 27509,
		617 => 27521,
		618 => 27532,
		619 => 27544,
		620 => 27556,
		621 => 27568,
		622 => 27579,
		623 => 27591,
		624 => 27603,
		625 => 27615,
		626 => 27626,
		627 => 27638,
		628 => 27649,
		629 => 27661,
		630 => 27673,
		631 => 27684,
		632 => 27696,
		633 => 27707,
		634 => 27719,
		635 => 27730,
		636 => 27742,
		637 => 27753,
		638 => 27764,
		639 => 27776,
		640 => 27787,
		641 => 27798,
		642 => 27810,
		643 => 27821,
		644 => 27832,
		645 => 27844,
		646 => 27855,
		647 => 27866,
		648 => 27877,
		649 => 27888,
		650 => 27900,
		651 => 27911,
		652 => 27922,
		653 => 27933,
		654 => 27944,
		655 => 27955,
		656 => 27966,
		657 => 27977,
		658 => 27988,
		659 => 27999,
		660 => 28010,
		661 => 28021,
		662 => 28032,
		663 => 28042,
		664 => 28053,
		665 => 28064,
		666 => 28075,
		667 => 28086,
		668 => 28097,
		669 => 28107,
		670 => 28118,
		671 => 28129,
		672 => 28139,
		673 => 28150,
		674 => 28161,
		675 => 28171,
		676 => 28182,
		677 => 28193,
		678 => 28203,
		679 => 28214,
		680 => 28224,
		681 => 28235,
		682 => 28245,
		683 => 28256,
		684 => 28266,
		685 => 28276,
		686 => 28287,
		687 => 28297,
		688 => 28308,
		689 => 28318,
		690 => 28328,
		691 => 28339,
		692 => 28349,
		693 => 28359,
		694 => 28369,
		695 => 28380,
		696 => 28390,
		697 => 28400,
		698 => 28410,
		699 => 28420,
		700 => 28430,
		701 => 28440,
		702 => 28450,
		703 => 28461,
		704 => 28471,
		705 => 28481,
		706 => 28491,
		707 => 28501,
		708 => 28511,
		709 => 28520,
		710 => 28530,
		711 => 28540,
		712 => 28550,
		713 => 28560,
		714 => 28570,
		715 => 28580,
		716 => 28589,
		717 => 28599,
		718 => 28609,
		719 => 28619,
		720 => 28628,
		721 => 28638,
		722 => 28648,
		723 => 28658,
		724 => 28667,
		725 => 28677,
		726 => 28686,
		727 => 28696,
		728 => 28706,
		729 => 28715,
		730 => 28725,
		731 => 28734,
		732 => 28744,
		733 => 28753,
		734 => 28763,
		735 => 28772,
		736 => 28781,
		737 => 28791,
		738 => 28800,
		739 => 28810,
		740 => 28819,
		741 => 28828,
		742 => 28837,
		743 => 28847,
		744 => 28856,
		745 => 28865,
		746 => 28874,
		747 => 28884,
		748 => 28893,
		749 => 28902,
		750 => 28911,
		751 => 28920,
		752 => 28929,
		753 => 28939,
		754 => 28948,
		755 => 28957,
		756 => 28966,
		757 => 28975,
		758 => 28984,
		759 => 28993,
		760 => 29002,
		761 => 29011,
		762 => 29020,
		763 => 29028,
		764 => 29037,
		765 => 29046,
		766 => 29055,
		767 => 29064,
		768 => 29073,
		769 => 29081,
		770 => 29090,
		771 => 29099,
		772 => 29108,
		773 => 29116,
		774 => 29125,
		775 => 29134,
		776 => 29143,
		777 => 29151,
		778 => 29160,
		779 => 29168,
		780 => 29177,
		781 => 29186,
		782 => 29194,
		783 => 29203,
		784 => 29211,
		785 => 29220,
		786 => 29228,
		787 => 29237,
		788 => 29245,
		789 => 29254,
		790 => 29262,
		791 => 29270,
		792 => 29279,
		793 => 29287,
		794 => 29295,
		795 => 29304,
		796 => 29312,
		797 => 29320,
		798 => 29329,
		799 => 29337,
		800 => 29345,
		801 => 29353,
		802 => 29362,
		803 => 29370,
		804 => 29378,
		805 => 29386,
		806 => 29394,
		807 => 29402,
		808 => 29410,
		809 => 29419,
		810 => 29427,
		811 => 29435,
		812 => 29443,
		813 => 29451,
		814 => 29459,
		815 => 29467,
		816 => 29475,
		817 => 29483,
		818 => 29491,
		819 => 29498,
		820 => 29506,
		821 => 29514,
		822 => 29522,
		823 => 29530,
		824 => 29538,
		825 => 29546,
		826 => 29553,
		827 => 29561,
		828 => 29569,
		829 => 29577,
		830 => 29584,
		831 => 29592,
		832 => 29600,
		833 => 29607,
		834 => 29615,
		835 => 29623,
		836 => 29630,
		837 => 29638,
		838 => 29646,
		839 => 29653,
		840 => 29661,
		841 => 29668,
		842 => 29676,
		843 => 29683,
		844 => 29691,
		845 => 29698,
		846 => 29706,
		847 => 29713,
		848 => 29721,
		849 => 29728,
		850 => 29735,
		851 => 29743,
		852 => 29750,
		853 => 29758,
		854 => 29765,
		855 => 29772,
		856 => 29780,
		857 => 29787,
		858 => 29794,
		859 => 29801,
		860 => 29809,
		861 => 29816,
		862 => 29823,
		863 => 29830,
		864 => 29837,
		865 => 29845,
		866 => 29852,
		867 => 29859,
		868 => 29866,
		869 => 29873,
		870 => 29880,
		871 => 29887,
		872 => 29894,
		873 => 29901,
		874 => 29908,
		875 => 29915,
		876 => 29922,
		877 => 29929,
		878 => 29936,
		879 => 29943,
		880 => 29950,
		881 => 29957,
		882 => 29964,
		883 => 29971,
		884 => 29978,
		885 => 29984,
		886 => 29991,
		887 => 29998,
		888 => 30005,
		889 => 30012,
		890 => 30018,
		891 => 30025,
		892 => 30032,
		893 => 30039,
		894 => 30045,
		895 => 30052,
		896 => 30059,
		897 => 30065,
		898 => 30072,
		899 => 30079,
		900 => 30085,
		901 => 30092,
		902 => 30098,
		903 => 30105,
		904 => 30112,
		905 => 30118,
		906 => 30125,
		907 => 30131,
		908 => 30138,
		909 => 30144,
		910 => 30151,
		911 => 30157,
		912 => 30164,
		913 => 30170,
		914 => 30176,
		915 => 30183,
		916 => 30189,
		917 => 30196,
		918 => 30202,
		919 => 30208,
		920 => 30215,
		921 => 30221,
		922 => 30227,
		923 => 30234,
		924 => 30240,
		925 => 30246,
		926 => 30252,
		927 => 30259,
		928 => 30265,
		929 => 30271,
		930 => 30277,
		931 => 30283,
		932 => 30289,
		933 => 30296,
		934 => 30302,
		935 => 30308,
		936 => 30314,
		937 => 30320,
		938 => 30326,
		939 => 30332,
		940 => 30338,
		941 => 30344,
		942 => 30350,
		943 => 30356,
		944 => 30362,
		945 => 30368,
		946 => 30374,
		947 => 30380,
		948 => 30386,
		949 => 30392,
		950 => 30398,
		951 => 30404,
		952 => 30410,
		953 => 30416,
		954 => 30421,
		955 => 30427,
		956 => 30433,
		957 => 30439,
		958 => 30445,
		959 => 30451,
		960 => 30456,
		961 => 30462,
		962 => 30468,
		963 => 30474,
		964 => 30479,
		965 => 30485,
		966 => 30491,
		967 => 30496,
		968 => 30502,
		969 => 30508,
		970 => 30513,
		971 => 30519,
		972 => 30525,
		973 => 30530,
		974 => 30536,
		975 => 30541,
		976 => 30547,
		977 => 30553,
		978 => 30558,
		979 => 30564,
		980 => 30569,
		981 => 30575,
		982 => 30580,
		983 => 30586,
		984 => 30591,
		985 => 30596,
		986 => 30602,
		987 => 30607,
		988 => 30613,
		989 => 30618,
		990 => 30624,
		991 => 30629,
		992 => 30634,
		993 => 30640,
		994 => 30645,
		995 => 30650,
		996 => 30656,
		997 => 30661,
		998 => 30666,
		999 => 30671,
		1000 => 30677,
		1001 => 30682,
		1002 => 30687,
		1003 => 30692,
		1004 => 30698,
		1005 => 30703,
		1006 => 30708,
		1007 => 30713,
		1008 => 30718,
		1009 => 30724,
		1010 => 30729,
		1011 => 30734,
		1012 => 30739,
		1013 => 30744,
		1014 => 30749,
		1015 => 30754,
		1016 => 30759,
		1017 => 30764,
		1018 => 30769,
		1019 => 30774,
		1020 => 30779,
		1021 => 30784,
		1022 => 30789,
		1023 => 30794,
		1024 => 30799,
		1025 => 30804,
		1026 => 30809,
		1027 => 30814,
		1028 => 30819,
		1029 => 30824,
		1030 => 30829,
		1031 => 30834,
		1032 => 30839,
		1033 => 30844,
		1034 => 30848,
		1035 => 30853,
		1036 => 30858,
		1037 => 30863,
		1038 => 30868,
		1039 => 30873,
		1040 => 30877,
		1041 => 30882,
		1042 => 30887,
		1043 => 30892,
		1044 => 30896,
		1045 => 30901,
		1046 => 30906,
		1047 => 30911,
		1048 => 30915,
		1049 => 30920,
		1050 => 30925,
		1051 => 30929,
		1052 => 30934,
		1053 => 30939,
		1054 => 30943,
		1055 => 30948,
		1056 => 30952,
		1057 => 30957,
		1058 => 30962,
		1059 => 30966,
		1060 => 30971,
		1061 => 30975,
		1062 => 30980,
		1063 => 30984,
		1064 => 30989,
		1065 => 30993,
		1066 => 30998,
		1067 => 31002,
		1068 => 31007,
		1069 => 31011,
		1070 => 31016,
		1071 => 31020,
		1072 => 31025,
		1073 => 31029,
		1074 => 31034,
		1075 => 31038,
		1076 => 31042,
		1077 => 31047,
		1078 => 31051,
		1079 => 31056,
		1080 => 31060,
		1081 => 31064,
		1082 => 31069,
		1083 => 31073,
		1084 => 31077,
		1085 => 31081,
		1086 => 31086,
		1087 => 31090,
		1088 => 31094,
		1089 => 31099,
		1090 => 31103,
		1091 => 31107,
		1092 => 31111,
		1093 => 31115,
		1094 => 31120,
		1095 => 31124,
		1096 => 31128,
		1097 => 31132,
		1098 => 31136,
		1099 => 31141,
		1100 => 31145,
		1101 => 31149,
		1102 => 31153,
		1103 => 31157,
		1104 => 31161,
		1105 => 31165,
		1106 => 31169,
		1107 => 31173,
		1108 => 31178,
		1109 => 31182,
		1110 => 31186,
		1111 => 31190,
		1112 => 31194,
		1113 => 31198,
		1114 => 31202,
		1115 => 31206,
		1116 => 31210,
		1117 => 31214,
		1118 => 31218,
		1119 => 31222,
		1120 => 31226,
		1121 => 31230,
		1122 => 31233,
		1123 => 31237,
		1124 => 31241,
		1125 => 31245,
		1126 => 31249,
		1127 => 31253,
		1128 => 31257,
		1129 => 31261,
		1130 => 31265,
		1131 => 31268,
		1132 => 31272,
		1133 => 31276,
		1134 => 31280,
		1135 => 31284,
		1136 => 31288,
		1137 => 31291,
		1138 => 31295,
		1139 => 31299,
		1140 => 31303,
		1141 => 31306,
		1142 => 31310,
		1143 => 31314,
		1144 => 31318,
		1145 => 31321,
		1146 => 31325,
		1147 => 31329,
		1148 => 31332,
		1149 => 31336,
		1150 => 31340,
		1151 => 31343,
		1152 => 31347,
		1153 => 31351,
		1154 => 31354,
		1155 => 31358,
		1156 => 31362,
		1157 => 31365,
		1158 => 31369,
		1159 => 31372,
		1160 => 31376,
		1161 => 31380,
		1162 => 31383,
		1163 => 31387,
		1164 => 31390,
		1165 => 31394,
		1166 => 31397,
		1167 => 31401,
		1168 => 31404,
		1169 => 31408,
		1170 => 31411,
		1171 => 31415,
		1172 => 31418,
		1173 => 31422,
		1174 => 31425,
		1175 => 31429,
		1176 => 31432,
		1177 => 31436,
		1178 => 31439,
		1179 => 31442,
		1180 => 31446,
		1181 => 31449,
		1182 => 31453,
		1183 => 31456,
		1184 => 31459,
		1185 => 31463,
		1186 => 31466,
		1187 => 31469,
		1188 => 31473,
		1189 => 31476,
		1190 => 31479,
		1191 => 31483,
		1192 => 31486,
		1193 => 31489,
		1194 => 31493,
		1195 => 31496,
		1196 => 31499,
		1197 => 31502,
		1198 => 31506,
		1199 => 31509,
		1200 => 31512,
		1201 => 31515,
		1202 => 31519,
		1203 => 31522,
		1204 => 31525,
		1205 => 31528,
		1206 => 31532,
		1207 => 31535,
		1208 => 31538,
		1209 => 31541,
		1210 => 31544,
		1211 => 31547,
		1212 => 31551,
		1213 => 31554,
		1214 => 31557,
		1215 => 31560,
		1216 => 31563,
		1217 => 31566,
		1218 => 31569,
		1219 => 31572,
		1220 => 31575,
		1221 => 31579,
		1222 => 31582,
		1223 => 31585,
		1224 => 31588,
		1225 => 31591,
		1226 => 31594,
		1227 => 31597,
		1228 => 31600,
		1229 => 31603,
		1230 => 31606,
		1231 => 31609,
		1232 => 31612,
		1233 => 31615,
		1234 => 31618,
		1235 => 31621,
		1236 => 31624,
		1237 => 31627,
		1238 => 31630,
		1239 => 31633,
		1240 => 31636,
		1241 => 31639,
		1242 => 31642,
		1243 => 31644,
		1244 => 31647,
		1245 => 31650,
		1246 => 31653,
		1247 => 31656,
		1248 => 31659,
		1249 => 31662,
		1250 => 31665,
		1251 => 31668,
		1252 => 31670,
		1253 => 31673,
		1254 => 31676,
		1255 => 31679,
		1256 => 31682,
		1257 => 31685,
		1258 => 31687,
		1259 => 31690,
		1260 => 31693,
		1261 => 31696,
		1262 => 31698,
		1263 => 31701,
		1264 => 31704,
		1265 => 31707,
		1266 => 31710,
		1267 => 31712,
		1268 => 31715,
		1269 => 31718,
		1270 => 31720,
		1271 => 31723,
		1272 => 31726,
		1273 => 31729,
		1274 => 31731,
		1275 => 31734,
		1276 => 31737,
		1277 => 31739,
		1278 => 31742,
		1279 => 31745,
		1280 => 31747,
		1281 => 31750,
		1282 => 31753,
		1283 => 31755,
		1284 => 31758,
		1285 => 31761,
		1286 => 31763,
		1287 => 31766,
		1288 => 31768,
		1289 => 31771,
		1290 => 31774,
		1291 => 31776,
		1292 => 31779,
		1293 => 31781,
		1294 => 31784,
		1295 => 31786,
		1296 => 31789,
		1297 => 31792,
		1298 => 31794,
		1299 => 31797,
		1300 => 31799,
		1301 => 31802,
		1302 => 31804,
		1303 => 31807,
		1304 => 31809,
		1305 => 31812,
		1306 => 31814,
		1307 => 31817,
		1308 => 31819,
		1309 => 31822,
		1310 => 31824,
		1311 => 31826,
		1312 => 31829,
		1313 => 31831,
		1314 => 31834,
		1315 => 31836,
		1316 => 31839,
		1317 => 31841,
		1318 => 31843,
		1319 => 31846,
		1320 => 31848,
		1321 => 31851,
		1322 => 31853,
		1323 => 31855,
		1324 => 31858,
		1325 => 31860,
		1326 => 31863,
		1327 => 31865,
		1328 => 31867,
		1329 => 31870,
		1330 => 31872,
		1331 => 31874,
		1332 => 31877,
		1333 => 31879,
		1334 => 31881,
		1335 => 31884,
		1336 => 31886,
		1337 => 31888,
		1338 => 31891,
		1339 => 31893,
		1340 => 31895,
		1341 => 31897,
		1342 => 31900,
		1343 => 31902,
		1344 => 31904,
		1345 => 31906,
		1346 => 31909,
		1347 => 31911,
		1348 => 31913,
		1349 => 31915,
		1350 => 31918,
		1351 => 31920,
		1352 => 31922,
		1353 => 31924,
		1354 => 31926,
		1355 => 31929,
		1356 => 31931,
		1357 => 31933,
		1358 => 31935,
		1359 => 31937,
		1360 => 31940,
		1361 => 31942,
		1362 => 31944,
		1363 => 31946,
		1364 => 31948,
		1365 => 31950,
		1366 => 31952,
		1367 => 31955,
		1368 => 31957,
		1369 => 31959,
		1370 => 31961,
		1371 => 31963,
		1372 => 31965,
		1373 => 31967,
		1374 => 31969,
		1375 => 31971,
		1376 => 31974,
		1377 => 31976,
		1378 => 31978,
		1379 => 31980,
		1380 => 31982,
		1381 => 31984,
		1382 => 31986,
		1383 => 31988,
		1384 => 31990,
		1385 => 31992,
		1386 => 31994,
		1387 => 31996,
		1388 => 31998,
		1389 => 32000,
		1390 => 32002,
		1391 => 32004,
		1392 => 32006,
		1393 => 32008,
		1394 => 32010,
		1395 => 32012,
		1396 => 32014,
		1397 => 32016,
		1398 => 32018,
		1399 => 32020,
		1400 => 32022,
		1401 => 32024,
		1402 => 32026,
		1403 => 32028,
		1404 => 32030,
		1405 => 32032,
		1406 => 32034,
		1407 => 32035,
		1408 => 32037,
		1409 => 32039,
		1410 => 32041,
		1411 => 32043,
		1412 => 32045,
		1413 => 32047,
		1414 => 32049,
		1415 => 32051,
		1416 => 32053,
		1417 => 32054,
		1418 => 32056,
		1419 => 32058,
		1420 => 32060,
		1421 => 32062,
		1422 => 32064,
		1423 => 32066,
		1424 => 32067,
		1425 => 32069,
		1426 => 32071,
		1427 => 32073,
		1428 => 32075,
		1429 => 32077,
		1430 => 32078,
		1431 => 32080,
		1432 => 32082,
		1433 => 32084,
		1434 => 32086,
		1435 => 32087,
		1436 => 32089,
		1437 => 32091,
		1438 => 32093,
		1439 => 32095,
		1440 => 32096,
		1441 => 32098,
		1442 => 32100,
		1443 => 32102,
		1444 => 32103,
		1445 => 32105,
		1446 => 32107,
		1447 => 32109,
		1448 => 32110,
		1449 => 32112,
		1450 => 32114,
		1451 => 32115,
		1452 => 32117,
		1453 => 32119,
		1454 => 32121,
		1455 => 32122,
		1456 => 32124,
		1457 => 32126,
		1458 => 32127,
		1459 => 32129,
		1460 => 32131,
		1461 => 32132,
		1462 => 32134,
		1463 => 32136,
		1464 => 32137,
		1465 => 32139,
		1466 => 32141,
		1467 => 32142,
		1468 => 32144,
		1469 => 32146,
		1470 => 32147,
		1471 => 32149,
		1472 => 32150,
		1473 => 32152,
		1474 => 32154,
		1475 => 32155,
		1476 => 32157,
		1477 => 32159,
		1478 => 32160,
		1479 => 32162,
		1480 => 32163,
		1481 => 32165,
		1482 => 32167,
		1483 => 32168,
		1484 => 32170,
		1485 => 32171,
		1486 => 32173,
		1487 => 32174,
		1488 => 32176,
		1489 => 32178,
		1490 => 32179,
		1491 => 32181,
		1492 => 32182,
		1493 => 32184,
		1494 => 32185,
		1495 => 32187,
		1496 => 32188,
		1497 => 32190,
		1498 => 32191,
		1499 => 32193,
		1500 => 32194,
		1501 => 32196,
		1502 => 32197,
		1503 => 32199,
		1504 => 32200,
		1505 => 32202,
		1506 => 32203,
		1507 => 32205,
		1508 => 32206,
		1509 => 32208,
		1510 => 32209,
		1511 => 32211,
		1512 => 32212,
		1513 => 32214,
		1514 => 32215,
		1515 => 32217,
		1516 => 32218,
		1517 => 32220,
		1518 => 32221,
		1519 => 32222,
		1520 => 32224,
		1521 => 32225,
		1522 => 32227,
		1523 => 32228,
		1524 => 32230,
		1525 => 32231,
		1526 => 32232,
		1527 => 32234,
		1528 => 32235,
		1529 => 32237,
		1530 => 32238,
		1531 => 32239,
		1532 => 32241,
		1533 => 32242,
		1534 => 32244,
		1535 => 32245,
		1536 => 32246,
		1537 => 32248,
		1538 => 32249,
		1539 => 32250,
		1540 => 32252,
		1541 => 32253,
		1542 => 32255,
		1543 => 32256,
		1544 => 32257,
		1545 => 32259,
		1546 => 32260,
		1547 => 32261,
		1548 => 32263,
		1549 => 32264,
		1550 => 32265,
		1551 => 32267,
		1552 => 32268,
		1553 => 32269,
		1554 => 32271,
		1555 => 32272,
		1556 => 32273,
		1557 => 32274,
		1558 => 32276,
		1559 => 32277,
		1560 => 32278,
		1561 => 32280,
		1562 => 32281,
		1563 => 32282,
		1564 => 32283,
		1565 => 32285,
		1566 => 32286,
		1567 => 32287,
		1568 => 32289,
		1569 => 32290,
		1570 => 32291,
		1571 => 32292,
		1572 => 32294,
		1573 => 32295,
		1574 => 32296,
		1575 => 32297,
		1576 => 32299,
		1577 => 32300,
		1578 => 32301,
		1579 => 32302,
		1580 => 32304,
		1581 => 32305,
		1582 => 32306,
		1583 => 32307,
		1584 => 32308,
		1585 => 32310,
		1586 => 32311,
		1587 => 32312,
		1588 => 32313,
		1589 => 32314,
		1590 => 32316,
		1591 => 32317,
		1592 => 32318,
		1593 => 32319,
		1594 => 32320,
		1595 => 32322,
		1596 => 32323,
		1597 => 32324,
		1598 => 32325,
		1599 => 32326,
		1600 => 32327,
		1601 => 32329,
		1602 => 32330,
		1603 => 32331,
		1604 => 32332,
		1605 => 32333,
		1606 => 32334,
		1607 => 32336,
		1608 => 32337,
		1609 => 32338,
		1610 => 32339,
		1611 => 32340,
		1612 => 32341,
		1613 => 32342,
		1614 => 32343,
		1615 => 32345,
		1616 => 32346,
		1617 => 32347,
		1618 => 32348,
		1619 => 32349,
		1620 => 32350,
		1621 => 32351,
		1622 => 32352,
		1623 => 32353,
		1624 => 32355,
		1625 => 32356,
		1626 => 32357,
		1627 => 32358,
		1628 => 32359,
		1629 => 32360,
		1630 => 32361,
		1631 => 32362,
		1632 => 32363,
		1633 => 32364,
		1634 => 32365,
		1635 => 32366,
		1636 => 32367,
		1637 => 32369,
		1638 => 32370,
		1639 => 32371,
		1640 => 32372,
		1641 => 32373,
		1642 => 32374,
		1643 => 32375,
		1644 => 32376,
		1645 => 32377,
		1646 => 32378,
		1647 => 32379,
		1648 => 32380,
		1649 => 32381,
		1650 => 32382,
		1651 => 32383,
		1652 => 32384,
		1653 => 32385,
		1654 => 32386,
		1655 => 32387,
		1656 => 32388,
		1657 => 32389,
		1658 => 32390,
		1659 => 32391,
		1660 => 32392,
		1661 => 32393,
		1662 => 32394,
		1663 => 32395,
		1664 => 32396,
		1665 => 32397,
		1666 => 32398,
		1667 => 32399,
		1668 => 32400,
		1669 => 32401,
		1670 => 32402,
		1671 => 32403,
		1672 => 32404,
		1673 => 32405,
		1674 => 32406,
		1675 => 32407,
		1676 => 32408,
		1677 => 32409,
		1678 => 32410,
		1679 => 32411,
		1680 => 32412,
		1681 => 32412,
		1682 => 32413,
		1683 => 32414,
		1684 => 32415,
		1685 => 32416,
		1686 => 32417,
		1687 => 32418,
		1688 => 32419,
		1689 => 32420,
		1690 => 32421,
		1691 => 32422,
		1692 => 32423,
		1693 => 32424,
		1694 => 32425,
		1695 => 32425,
		1696 => 32426,
		1697 => 32427,
		1698 => 32428,
		1699 => 32429,
		1700 => 32430,
		1701 => 32431,
		1702 => 32432,
		1703 => 32433,
		1704 => 32433,
		1705 => 32434,
		1706 => 32435,
		1707 => 32436,
		1708 => 32437,
		1709 => 32438,
		1710 => 32439,
		1711 => 32440,
		1712 => 32441,
		1713 => 32441,
		1714 => 32442,
		1715 => 32443,
		1716 => 32444,
		1717 => 32445,
		1718 => 32446,
		1719 => 32447,
		1720 => 32447,
		1721 => 32448,
		1722 => 32449,
		1723 => 32450,
		1724 => 32451,
		1725 => 32452,
		1726 => 32452,
		1727 => 32453,
		1728 => 32454,
		1729 => 32455,
		1730 => 32456,
		1731 => 32457,
		1732 => 32457,
		1733 => 32458,
		1734 => 32459,
		1735 => 32460,
		1736 => 32461,
		1737 => 32462,
		1738 => 32462,
		1739 => 32463,
		1740 => 32464,
		1741 => 32465,
		1742 => 32466,
		1743 => 32466,
		1744 => 32467,
		1745 => 32468,
		1746 => 32469,
		1747 => 32470,
		1748 => 32470,
		1749 => 32471,
		1750 => 32472,
		1751 => 32473,
		1752 => 32473,
		1753 => 32474,
		1754 => 32475,
		1755 => 32476,
		1756 => 32477,
		1757 => 32477,
		1758 => 32478,
		1759 => 32479,
		1760 => 32480,
		1761 => 32480,
		1762 => 32481,
		1763 => 32482,
		1764 => 32483,
		1765 => 32483,
		1766 => 32484,
		1767 => 32485,
		1768 => 32486,
		1769 => 32486,
		1770 => 32487,
		1771 => 32488,
		1772 => 32489,
		1773 => 32489,
		1774 => 32490,
		1775 => 32491,
		1776 => 32492,
		1777 => 32492,
		1778 => 32493,
		1779 => 32494,
		1780 => 32495,
		1781 => 32495,
		1782 => 32496,
		1783 => 32497,
		1784 => 32497,
		1785 => 32498,
		1786 => 32499,
		1787 => 32500,
		1788 => 32500,
		1789 => 32501,
		1790 => 32502,
		1791 => 32502,
		1792 => 32503,
		1793 => 32504,
		1794 => 32505,
		1795 => 32505,
		1796 => 32506,
		1797 => 32507,
		1798 => 32507,
		1799 => 32508,
		1800 => 32509,
		1801 => 32509,
		1802 => 32510,
		1803 => 32511,
		1804 => 32511,
		1805 => 32512,
		1806 => 32513,
		1807 => 32513,
		1808 => 32514,
		1809 => 32515,
		1810 => 32515,
		1811 => 32516,
		1812 => 32517,
		1813 => 32518,
		1814 => 32518,
		1815 => 32519,
		1816 => 32519,
		1817 => 32520,
		1818 => 32521,
		1819 => 32521,
		1820 => 32522,
		1821 => 32523,
		1822 => 32523,
		1823 => 32524,
		1824 => 32525,
		1825 => 32525,
		1826 => 32526,
		1827 => 32527,
		1828 => 32527,
		1829 => 32528,
		1830 => 32529,
		1831 => 32529,
		1832 => 32530,
		1833 => 32530,
		1834 => 32531,
		1835 => 32532,
		1836 => 32532,
		1837 => 32533,
		1838 => 32534,
		1839 => 32534,
		1840 => 32535,
		1841 => 32535,
		1842 => 32536,
		1843 => 32537,
		1844 => 32537,
		1845 => 32538,
		1846 => 32539,
		1847 => 32539,
		1848 => 32540,
		1849 => 32540,
		1850 => 32541,
		1851 => 32542,
		1852 => 32542,
		1853 => 32543,
		1854 => 32543,
		1855 => 32544,
		1856 => 32545,
		1857 => 32545,
		1858 => 32546,
		1859 => 32546,
		1860 => 32547,
		1861 => 32547,
		1862 => 32548,
		1863 => 32549,
		1864 => 32549,
		1865 => 32550,
		1866 => 32550,
		1867 => 32551,
		1868 => 32552,
		1869 => 32552,
		1870 => 32553,
		1871 => 32553,
		1872 => 32554,
		1873 => 32554,
		1874 => 32555,
		1875 => 32556,
		1876 => 32556,
		1877 => 32557,
		1878 => 32557,
		1879 => 32558,
		1880 => 32558,
		1881 => 32559,
		1882 => 32559,
		1883 => 32560,
		1884 => 32561,
		1885 => 32561,
		1886 => 32562,
		1887 => 32562,
		1888 => 32563,
		1889 => 32563,
		1890 => 32564,
		1891 => 32564,
		1892 => 32565,
		1893 => 32565,
		1894 => 32566,
		1895 => 32567,
		1896 => 32567,
		1897 => 32568,
		1898 => 32568,
		1899 => 32569,
		1900 => 32569,
		1901 => 32570,
		1902 => 32570,
		1903 => 32571,
		1904 => 32571,
		1905 => 32572,
		1906 => 32572,
		1907 => 32573,
		1908 => 32573,
		1909 => 32574,
		1910 => 32574,
		1911 => 32575,
		1912 => 32575,
		1913 => 32576,
		1914 => 32576,
		1915 => 32577,
		1916 => 32577,
		1917 => 32578,
		1918 => 32578,
		1919 => 32579,
		1920 => 32579,
		1921 => 32580,
		1922 => 32580,
		1923 => 32581,
		1924 => 32581,
		1925 => 32582,
		1926 => 32582,
		1927 => 32583,
		1928 => 32583,
		1929 => 32584,
		1930 => 32584,
		1931 => 32585,
		1932 => 32585,
		1933 => 32586,
		1934 => 32586,
		1935 => 32587,
		1936 => 32587,
		1937 => 32588,
		1938 => 32588,
		1939 => 32589,
		1940 => 32589,
		1941 => 32590,
		1942 => 32590,
		1943 => 32591,
		1944 => 32591,
		1945 => 32592,
		1946 => 32592,
		1947 => 32593,
		1948 => 32593,
		1949 => 32593,
		1950 => 32594,
		1951 => 32594,
		1952 => 32595,
		1953 => 32595,
		1954 => 32596,
		1955 => 32596,
		1956 => 32597,
		1957 => 32597,
		1958 => 32598,
		1959 => 32598,
		1960 => 32598,
		1961 => 32599,
		1962 => 32599,
		1963 => 32600,
		1964 => 32600,
		1965 => 32601,
		1966 => 32601,
		1967 => 32602,
		1968 => 32602,
		1969 => 32602,
		1970 => 32603,
		1971 => 32603,
		1972 => 32604,
		1973 => 32604,
		1974 => 32605,
		1975 => 32605,
		1976 => 32606,
		1977 => 32606,
		1978 => 32606,
		1979 => 32607,
		1980 => 32607,
		1981 => 32608,
		1982 => 32608,
		1983 => 32609,
		1984 => 32609,
		1985 => 32609,
		1986 => 32610,
		1987 => 32610,
		1988 => 32611,
		1989 => 32611,
		1990 => 32611,
		1991 => 32612,
		1992 => 32612,
		1993 => 32613,
		1994 => 32613,
		1995 => 32614,
		1996 => 32614,
		1997 => 32614,
		1998 => 32615,
		1999 => 32615,
		2000 => 32616,
		2001 => 32616,
		2002 => 32616,
		2003 => 32617,
		2004 => 32617,
		2005 => 32618,
		2006 => 32618,
		2007 => 32618,
		2008 => 32619,
		2009 => 32619,
		2010 => 32620,
		2011 => 32620,
		2012 => 32620,
		2013 => 32621,
		2014 => 32621,
		2015 => 32622,
		2016 => 32622,
		2017 => 32622,
		2018 => 32623,
		2019 => 32623,
		2020 => 32623,
		2021 => 32624,
		2022 => 32624,
		2023 => 32625,
		2024 => 32625,
		2025 => 32625,
		2026 => 32626,
		2027 => 32626,
		2028 => 32626,
		2029 => 32627,
		2030 => 32627,
		2031 => 32628,
		2032 => 32628,
		2033 => 32628,
		2034 => 32629,
		2035 => 32629,
		2036 => 32629,
		2037 => 32630,
		2038 => 32630,
		2039 => 32631,
		2040 => 32631,
		2041 => 32631,
		2042 => 32632,
		2043 => 32632,
		2044 => 32632,
		2045 => 32633,
		2046 => 32633,
		2047 => 32633,
		2048 => 32634,
		2049 => 32634,
		2050 => 32635,
		2051 => 32635,
		2052 => 32635,
		2053 => 32636,
		2054 => 32636,
		2055 => 32636,
		2056 => 32637,
		2057 => 32637,
		2058 => 32637,
		2059 => 32638,
		2060 => 32638,
		2061 => 32638,
		2062 => 32639,
		2063 => 32639,
		2064 => 32639,
		2065 => 32640,
		2066 => 32640,
		2067 => 32640,
		2068 => 32641,
		2069 => 32641,
		2070 => 32641,
		2071 => 32642,
		2072 => 32642,
		2073 => 32642,
		2074 => 32643,
		2075 => 32643,
		2076 => 32643,
		2077 => 32644,
		2078 => 32644,
		2079 => 32644,
		2080 => 32645,
		2081 => 32645,
		2082 => 32645,
		2083 => 32646,
		2084 => 32646,
		2085 => 32646,
		2086 => 32647,
		2087 => 32647,
		2088 => 32647,
		2089 => 32648,
		2090 => 32648,
		2091 => 32648,
		2092 => 32649,
		2093 => 32649,
		2094 => 32649,
		2095 => 32650,
		2096 => 32650,
		2097 => 32650,
		2098 => 32650,
		2099 => 32651,
		2100 => 32651,
		2101 => 32651,
		2102 => 32652,
		2103 => 32652,
		2104 => 32652,
		2105 => 32653,
		2106 => 32653,
		2107 => 32653,
		2108 => 32654,
		2109 => 32654,
		2110 => 32654,
		2111 => 32654,
		2112 => 32655,
		2113 => 32655,
		2114 => 32655,
		2115 => 32656,
		2116 => 32656,
		2117 => 32656,
		2118 => 32657,
		2119 => 32657,
		2120 => 32657,
		2121 => 32657,
		2122 => 32658,
		2123 => 32658,
		2124 => 32658,
		2125 => 32659,
		2126 => 32659,
		2127 => 32659,
		2128 => 32659,
		2129 => 32660,
		2130 => 32660,
		2131 => 32660,
		2132 => 32661,
		2133 => 32661,
		2134 => 32661,
		2135 => 32661,
		2136 => 32662,
		2137 => 32662,
		2138 => 32662,
		2139 => 32663,
		2140 => 32663,
		2141 => 32663,
		2142 => 32663,
		2143 => 32664,
		2144 => 32664,
		2145 => 32664,
		2146 => 32665,
		2147 => 32665,
		2148 => 32665,
		2149 => 32665,
		2150 => 32666,
		2151 => 32666,
		2152 => 32666,
		2153 => 32666,
		2154 => 32667,
		2155 => 32667,
		2156 => 32667,
		2157 => 32668,
		2158 => 32668,
		2159 => 32668,
		2160 => 32668,
		2161 => 32669,
		2162 => 32669,
		2163 => 32669,
		2164 => 32669,
		2165 => 32670,
		2166 => 32670,
		2167 => 32670,
		2168 => 32670,
		2169 => 32671,
		2170 => 32671,
		2171 => 32671,
		2172 => 32671,
		2173 => 32672,
		2174 => 32672,
		2175 => 32672,
		2176 => 32672,
		2177 => 32673,
		2178 => 32673,
		2179 => 32673,
		2180 => 32673,
		2181 => 32674,
		2182 => 32674,
		2183 => 32674,
		2184 => 32674,
		2185 => 32675,
		2186 => 32675,
		2187 => 32675,
		2188 => 32675,
		2189 => 32676,
		2190 => 32676,
		2191 => 32676,
		2192 => 32676,
		2193 => 32677,
		2194 => 32677,
		2195 => 32677,
		2196 => 32677,
		2197 => 32678,
		2198 => 32678,
		2199 => 32678,
		2200 => 32678,
		2201 => 32679,
		2202 => 32679,
		2203 => 32679,
		2204 => 32679,
		2205 => 32680,
		2206 => 32680,
		2207 => 32680,
		2208 => 32680,
		2209 => 32680,
		2210 => 32681,
		2211 => 32681,
		2212 => 32681,
		2213 => 32681,
		2214 => 32682,
		2215 => 32682,
		2216 => 32682,
		2217 => 32682,
		2218 => 32683,
		2219 => 32683,
		2220 => 32683,
		2221 => 32683,
		2222 => 32683,
		2223 => 32684,
		2224 => 32684,
		2225 => 32684,
		2226 => 32684,
		2227 => 32685,
		2228 => 32685,
		2229 => 32685,
		2230 => 32685,
		2231 => 32685,
		2232 => 32686,
		2233 => 32686,
		2234 => 32686,
		2235 => 32686,
		2236 => 32686,
		2237 => 32687,
		2238 => 32687,
		2239 => 32687,
		2240 => 32687,
		2241 => 32688,
		2242 => 32688,
		2243 => 32688,
		2244 => 32688,
		2245 => 32688,
		2246 => 32689,
		2247 => 32689,
		2248 => 32689,
		2249 => 32689,
		2250 => 32689,
		2251 => 32690,
		2252 => 32690,
		2253 => 32690,
		2254 => 32690,
		2255 => 32690,
		2256 => 32691,
		2257 => 32691,
		2258 => 32691,
		2259 => 32691,
		2260 => 32692,
		2261 => 32692,
		2262 => 32692,
		2263 => 32692,
		2264 => 32692,
		2265 => 32693,
		2266 => 32693,
		2267 => 32693,
		2268 => 32693,
		2269 => 32693,
		2270 => 32694,
		2271 => 32694,
		2272 => 32694,
		2273 => 32694,
		2274 => 32694,
		2275 => 32694,
		2276 => 32695,
		2277 => 32695,
		2278 => 32695,
		2279 => 32695,
		2280 => 32695,
		2281 => 32696,
		2282 => 32696,
		2283 => 32696,
		2284 => 32696,
		2285 => 32696,
		2286 => 32697,
		2287 => 32697,
		2288 => 32697,
		2289 => 32697,
		2290 => 32697,
		2291 => 32698,
		2292 => 32698,
		2293 => 32698,
		2294 => 32698,
		2295 => 32698,
		2296 => 32698,
		2297 => 32699,
		2298 => 32699,
		2299 => 32699,
		2300 => 32699,
		2301 => 32699,
		2302 => 32700,
		2303 => 32700,
		2304 => 32700,
		2305 => 32700,
		2306 => 32700,
		2307 => 32700,
		2308 => 32701,
		2309 => 32701,
		2310 => 32701,
		2311 => 32701,
		2312 => 32701,
		2313 => 32702,
		2314 => 32702,
		2315 => 32702,
		2316 => 32702,
		2317 => 32702,
		2318 => 32702,
		2319 => 32703,
		2320 => 32703,
		2321 => 32703,
		2322 => 32703,
		2323 => 32703,
		2324 => 32703,
		2325 => 32704,
		2326 => 32704,
		2327 => 32704,
		2328 => 32704,
		2329 => 32704,
		2330 => 32704,
		2331 => 32705,
		2332 => 32705,
		2333 => 32705,
		2334 => 32705,
		2335 => 32705,
		2336 => 32705,
		2337 => 32706,
		2338 => 32706,
		2339 => 32706,
		2340 => 32706,
		2341 => 32706,
		2342 => 32706,
		2343 => 32707,
		2344 => 32707,
		2345 => 32707,
		2346 => 32707,
		2347 => 32707,
		2348 => 32707,
		2349 => 32708,
		2350 => 32708,
		2351 => 32708,
		2352 => 32708,
		2353 => 32708,
		2354 => 32708,
		2355 => 32708,
		2356 => 32709,
		2357 => 32709,
		2358 => 32709,
		2359 => 32709,
		2360 => 32709,
		2361 => 32709,
		2362 => 32710,
		2363 => 32710,
		2364 => 32710,
		2365 => 32710,
		2366 => 32710,
		2367 => 32710,
		2368 => 32710,
		2369 => 32711,
		2370 => 32711,
		2371 => 32711,
		2372 => 32711,
		2373 => 32711,
		2374 => 32711,
		2375 => 32712,
		2376 => 32712,
		2377 => 32712,
		2378 => 32712,
		2379 => 32712,
		2380 => 32712,
		2381 => 32712,
		2382 => 32713,
		2383 => 32713,
		2384 => 32713,
		2385 => 32713,
		2386 => 32713,
		2387 => 32713,
		2388 => 32713,
		2389 => 32714,
		2390 => 32714,
		2391 => 32714,
		2392 => 32714,
		2393 => 32714,
		2394 => 32714,
		2395 => 32714,
		2396 => 32715,
		2397 => 32715,
		2398 => 32715,
		2399 => 32715,
		2400 => 32715,
		2401 => 32715,
		2402 => 32715,
		2403 => 32716,
		2404 => 32716,
		2405 => 32716,
		2406 => 32716,
		2407 => 32716,
		2408 => 32716,
		2409 => 32716,
		2410 => 32717,
		2411 => 32717,
		2412 => 32717,
		2413 => 32717,
		2414 => 32717,
		2415 => 32717,
		2416 => 32717,
		2417 => 32717,
		2418 => 32718,
		2419 => 32718,
		2420 => 32718,
		2421 => 32718,
		2422 => 32718,
		2423 => 32718,
		2424 => 32718,
		2425 => 32718,
		2426 => 32719,
		2427 => 32719,
		2428 => 32719,
		2429 => 32719,
		2430 => 32719,
		2431 => 32719,
		2432 => 32719,
		2433 => 32720,
		2434 => 32720,
		2435 => 32720,
		2436 => 32720,
		2437 => 32720,
		2438 => 32720,
		2439 => 32720,
		2440 => 32720,
		2441 => 32721,
		2442 => 32721,
		2443 => 32721,
		2444 => 32721,
		2445 => 32721,
		2446 => 32721,
		2447 => 32721,
		2448 => 32721,
		2449 => 32722,
		2450 => 32722,
		2451 => 32722,
		2452 => 32722,
		2453 => 32722,
		2454 => 32722,
		2455 => 32722,
		2456 => 32722,
		2457 => 32722,
		2458 => 32723,
		2459 => 32723,
		2460 => 32723,
		2461 => 32723,
		2462 => 32723,
		2463 => 32723,
		2464 => 32723,
		2465 => 32723,
		2466 => 32724,
		2467 => 32724,
		2468 => 32724,
		2469 => 32724,
		2470 => 32724,
		2471 => 32724,
		2472 => 32724,
		2473 => 32724,
		2474 => 32724,
		2475 => 32725,
		2476 => 32725,
		2477 => 32725,
		2478 => 32725,
		2479 => 32725,
		2480 => 32725,
		2481 => 32725,
		2482 => 32725,
		2483 => 32725,
		2484 => 32726,
		2485 => 32726,
		2486 => 32726,
		2487 => 32726,
		2488 => 32726,
		2489 => 32726,
		2490 => 32726,
		2491 => 32726,
		2492 => 32726,
		2493 => 32727,
		2494 => 32727,
		2495 => 32727,
		2496 => 32727,
		2497 => 32727,
		2498 => 32727,
		2499 => 32727,
		2500 => 32727,
		2501 => 32727,
		2502 => 32728,
		2503 => 32728,
		2504 => 32728,
		2505 => 32728,
		2506 => 32728,
		2507 => 32728,
		2508 => 32728,
		2509 => 32728,
		2510 => 32728,
		2511 => 32728,
		2512 => 32729,
		2513 => 32729,
		2514 => 32729,
		2515 => 32729,
		2516 => 32729,
		2517 => 32729,
		2518 => 32729,
		2519 => 32729,
		2520 => 32729,
		2521 => 32730,
		2522 => 32730,
		2523 => 32730,
		2524 => 32730,
		2525 => 32730,
		2526 => 32730,
		2527 => 32730,
		2528 => 32730,
		2529 => 32730,
		2530 => 32730,
		2531 => 32731,
		2532 => 32731,
		2533 => 32731,
		2534 => 32731,
		2535 => 32731,
		2536 => 32731,
		2537 => 32731,
		2538 => 32731,
		2539 => 32731,
		2540 => 32731,
		2541 => 32731,
		2542 => 32732,
		2543 => 32732,
		2544 => 32732,
		2545 => 32732,
		2546 => 32732,
		2547 => 32732,
		2548 => 32732,
		2549 => 32732,
		2550 => 32732,
		2551 => 32732,
		2552 => 32733,
		2553 => 32733,
		2554 => 32733,
		2555 => 32733,
		2556 => 32733,
		2557 => 32733,
		2558 => 32733,
		2559 => 32733,
		2560 => 32733,
		2561 => 32733,
		2562 => 32733,
		2563 => 32734,
		2564 => 32734,
		2565 => 32734,
		2566 => 32734,
		2567 => 32734,
		2568 => 32734,
		2569 => 32734,
		2570 => 32734,
		2571 => 32734,
		2572 => 32734,
		2573 => 32734,
		2574 => 32734,
		2575 => 32735,
		2576 => 32735,
		2577 => 32735,
		2578 => 32735,
		2579 => 32735,
		2580 => 32735,
		2581 => 32735,
		2582 => 32735,
		2583 => 32735,
		2584 => 32735,
		2585 => 32735,
		2586 => 32736,
		2587 => 32736,
		2588 => 32736,
		2589 => 32736,
		2590 => 32736,
		2591 => 32736,
		2592 => 32736,
		2593 => 32736,
		2594 => 32736,
		2595 => 32736,
		2596 => 32736,
		2597 => 32736,
		2598 => 32737,
		2599 => 32737,
		2600 => 32737,
		2601 => 32737,
		2602 => 32737,
		2603 => 32737,
		2604 => 32737,
		2605 => 32737,
		2606 => 32737,
		2607 => 32737,
		2608 => 32737,
		2609 => 32737,
		2610 => 32737,
		2611 => 32738,
		2612 => 32738,
		2613 => 32738,
		2614 => 32738,
		2615 => 32738,
		2616 => 32738,
		2617 => 32738,
		2618 => 32738,
		2619 => 32738,
		2620 => 32738,
		2621 => 32738,
		2622 => 32738,
		2623 => 32738,
		2624 => 32739,
		2625 => 32739,
		2626 => 32739,
		2627 => 32739,
		2628 => 32739,
		2629 => 32739,
		2630 => 32739,
		2631 => 32739,
		2632 => 32739,
		2633 => 32739,
		2634 => 32739,
		2635 => 32739,
		2636 => 32739,
		2637 => 32740,
		2638 => 32740,
		2639 => 32740,
		2640 => 32740,
		2641 => 32740,
		2642 => 32740,
		2643 => 32740,
		2644 => 32740,
		2645 => 32740,
		2646 => 32740,
		2647 => 32740,
		2648 => 32740,
		2649 => 32740,
		2650 => 32740,
		2651 => 32741,
		2652 => 32741,
		2653 => 32741,
		2654 => 32741,
		2655 => 32741,
		2656 => 32741,
		2657 => 32741,
		2658 => 32741,
		2659 => 32741,
		2660 => 32741,
		2661 => 32741,
		2662 => 32741,
		2663 => 32741,
		2664 => 32741,
		2665 => 32742,
		2666 => 32742,
		2667 => 32742,
		2668 => 32742,
		2669 => 32742,
		2670 => 32742,
		2671 => 32742,
		2672 => 32742,
		2673 => 32742,
		2674 => 32742,
		2675 => 32742,
		2676 => 32742,
		2677 => 32742,
		2678 => 32742,
		2679 => 32742,
		2680 => 32743,
		2681 => 32743,
		2682 => 32743,
		2683 => 32743,
		2684 => 32743,
		2685 => 32743,
		2686 => 32743,
		2687 => 32743,
		2688 => 32743,
		2689 => 32743,
		2690 => 32743,
		2691 => 32743,
		2692 => 32743,
		2693 => 32743,
		2694 => 32743,
		2695 => 32743,
		2696 => 32744,
		2697 => 32744,
		2698 => 32744,
		2699 => 32744,
		2700 => 32744,
		2701 => 32744,
		2702 => 32744,
		2703 => 32744,
		2704 => 32744,
		2705 => 32744,
		2706 => 32744,
		2707 => 32744,
		2708 => 32744,
		2709 => 32744,
		2710 => 32744,
		2711 => 32744,
		2712 => 32745,
		2713 => 32745,
		2714 => 32745,
		2715 => 32745,
		2716 => 32745,
		2717 => 32745,
		2718 => 32745,
		2719 => 32745,
		2720 => 32745,
		2721 => 32745,
		2722 => 32745,
		2723 => 32745,
		2724 => 32745,
		2725 => 32745,
		2726 => 32745,
		2727 => 32745,
		2728 => 32745,
		2729 => 32746,
		2730 => 32746,
		2731 => 32746,
		2732 => 32746,
		2733 => 32746,
		2734 => 32746,
		2735 => 32746,
		2736 => 32746,
		2737 => 32746,
		2738 => 32746,
		2739 => 32746,
		2740 => 32746,
		2741 => 32746,
		2742 => 32746,
		2743 => 32746,
		2744 => 32746,
		2745 => 32746,
		2746 => 32747,
		2747 => 32747,
		2748 => 32747,
		2749 => 32747,
		2750 => 32747,
		2751 => 32747,
		2752 => 32747,
		2753 => 32747,
		2754 => 32747,
		2755 => 32747,
		2756 => 32747,
		2757 => 32747,
		2758 => 32747,
		2759 => 32747,
		2760 => 32747,
		2761 => 32747,
		2762 => 32747,
		2763 => 32747,
		2764 => 32747,
		2765 => 32748,
		2766 => 32748,
		2767 => 32748,
		2768 => 32748,
		2769 => 32748,
		2770 => 32748,
		2771 => 32748,
		2772 => 32748,
		2773 => 32748,
		2774 => 32748,
		2775 => 32748,
		2776 => 32748,
		2777 => 32748,
		2778 => 32748,
		2779 => 32748,
		2780 => 32748,
		2781 => 32748,
		2782 => 32748,
		2783 => 32748,
		2784 => 32748,
		2785 => 32749,
		2786 => 32749,
		2787 => 32749,
		2788 => 32749,
		2789 => 32749,
		2790 => 32749,
		2791 => 32749,
		2792 => 32749,
		2793 => 32749,
		2794 => 32749,
		2795 => 32749,
		2796 => 32749,
		2797 => 32749,
		2798 => 32749,
		2799 => 32749,
		2800 => 32749,
		2801 => 32749,
		2802 => 32749,
		2803 => 32749,
		2804 => 32749,
		2805 => 32750,
		2806 => 32750,
		2807 => 32750,
		2808 => 32750,
		2809 => 32750,
		2810 => 32750,
		2811 => 32750,
		2812 => 32750,
		2813 => 32750,
		2814 => 32750,
		2815 => 32750,
		2816 => 32750,
		2817 => 32750,
		2818 => 32750,
		2819 => 32750,
		2820 => 32750,
		2821 => 32750,
		2822 => 32750,
		2823 => 32750,
		2824 => 32750,
		2825 => 32750,
		2826 => 32750,
		2827 => 32751,
		2828 => 32751,
		2829 => 32751,
		2830 => 32751,
		2831 => 32751,
		2832 => 32751,
		2833 => 32751,
		2834 => 32751,
		2835 => 32751,
		2836 => 32751,
		2837 => 32751,
		2838 => 32751,
		2839 => 32751,
		2840 => 32751,
		2841 => 32751,
		2842 => 32751,
		2843 => 32751,
		2844 => 32751,
		2845 => 32751,
		2846 => 32751,
		2847 => 32751,
		2848 => 32751,
		2849 => 32751,
		2850 => 32751,
		2851 => 32752,
		2852 => 32752,
		2853 => 32752,
		2854 => 32752,
		2855 => 32752,
		2856 => 32752,
		2857 => 32752,
		2858 => 32752,
		2859 => 32752,
		2860 => 32752,
		2861 => 32752,
		2862 => 32752,
		2863 => 32752,
		2864 => 32752,
		2865 => 32752,
		2866 => 32752,
		2867 => 32752,
		2868 => 32752,
		2869 => 32752,
		2870 => 32752,
		2871 => 32752,
		2872 => 32752,
		2873 => 32752,
		2874 => 32752,
		2875 => 32753,
		2876 => 32753,
		2877 => 32753,
		2878 => 32753,
		2879 => 32753,
		2880 => 32753,
		2881 => 32753,
		2882 => 32753,
		2883 => 32753,
		2884 => 32753,
		2885 => 32753,
		2886 => 32753,
		2887 => 32753,
		2888 => 32753,
		2889 => 32753,
		2890 => 32753,
		2891 => 32753,
		2892 => 32753,
		2893 => 32753,
		2894 => 32753,
		2895 => 32753,
		2896 => 32753,
		2897 => 32753,
		2898 => 32753,
		2899 => 32753,
		2900 => 32753,
		2901 => 32753,
		2902 => 32754,
		2903 => 32754,
		2904 => 32754,
		2905 => 32754,
		2906 => 32754,
		2907 => 32754,
		2908 => 32754,
		2909 => 32754,
		2910 => 32754,
		2911 => 32754,
		2912 => 32754,
		2913 => 32754,
		2914 => 32754,
		2915 => 32754,
		2916 => 32754,
		2917 => 32754,
		2918 => 32754,
		2919 => 32754,
		2920 => 32754,
		2921 => 32754,
		2922 => 32754,
		2923 => 32754,
		2924 => 32754,
		2925 => 32754,
		2926 => 32754,
		2927 => 32754,
		2928 => 32754,
		2929 => 32754,
		2930 => 32754,
		2931 => 32755,
		2932 => 32755,
		2933 => 32755,
		2934 => 32755,
		2935 => 32755,
		2936 => 32755,
		2937 => 32755,
		2938 => 32755,
		2939 => 32755,
		2940 => 32755,
		2941 => 32755,
		2942 => 32755,
		2943 => 32755,
		2944 => 32755,
		2945 => 32755,
		2946 => 32755,
		2947 => 32755,
		2948 => 32755,
		2949 => 32755,
		2950 => 32755,
		2951 => 32755,
		2952 => 32755,
		2953 => 32755,
		2954 => 32755,
		2955 => 32755,
		2956 => 32755,
		2957 => 32755,
		2958 => 32755,
		2959 => 32755,
		2960 => 32755,
		2961 => 32755,
		2962 => 32756,
		2963 => 32756,
		2964 => 32756,
		2965 => 32756,
		2966 => 32756,
		2967 => 32756,
		2968 => 32756,
		2969 => 32756,
		2970 => 32756,
		2971 => 32756,
		2972 => 32756,
		2973 => 32756,
		2974 => 32756,
		2975 => 32756,
		2976 => 32756,
		2977 => 32756,
		2978 => 32756,
		2979 => 32756,
		2980 => 32756,
		2981 => 32756,
		2982 => 32756,
		2983 => 32756,
		2984 => 32756,
		2985 => 32756,
		2986 => 32756,
		2987 => 32756,
		2988 => 32756,
		2989 => 32756,
		2990 => 32756,
		2991 => 32756,
		2992 => 32756,
		2993 => 32756,
		2994 => 32756,
		2995 => 32756,
		2996 => 32757,
		2997 => 32757,
		2998 => 32757,
		2999 => 32757,
		3000 => 32757,
		3001 => 32757,
		3002 => 32757,
		3003 => 32757,
		3004 => 32757,
		3005 => 32757,
		3006 => 32757,
		3007 => 32757,
		3008 => 32757,
		3009 => 32757,
		3010 => 32757,
		3011 => 32757,
		3012 => 32757,
		3013 => 32757,
		3014 => 32757,
		3015 => 32757,
		3016 => 32757,
		3017 => 32757,
		3018 => 32757,
		3019 => 32757,
		3020 => 32757,
		3021 => 32757,
		3022 => 32757,
		3023 => 32757,
		3024 => 32757,
		3025 => 32757,
		3026 => 32757,
		3027 => 32757,
		3028 => 32757,
		3029 => 32757,
		3030 => 32757,
		3031 => 32757,
		3032 => 32757,
		3033 => 32758,
		3034 => 32758,
		3035 => 32758,
		3036 => 32758,
		3037 => 32758,
		3038 => 32758,
		3039 => 32758,
		3040 => 32758,
		3041 => 32758,
		3042 => 32758,
		3043 => 32758,
		3044 => 32758,
		3045 => 32758,
		3046 => 32758,
		3047 => 32758,
		3048 => 32758,
		3049 => 32758,
		3050 => 32758,
		3051 => 32758,
		3052 => 32758,
		3053 => 32758,
		3054 => 32758,
		3055 => 32758,
		3056 => 32758,
		3057 => 32758,
		3058 => 32758,
		3059 => 32758,
		3060 => 32758,
		3061 => 32758,
		3062 => 32758,
		3063 => 32758,
		3064 => 32758,
		3065 => 32758,
		3066 => 32758,
		3067 => 32758,
		3068 => 32758,
		3069 => 32758,
		3070 => 32758,
		3071 => 32758,
		3072 => 32758,
		3073 => 32758,
		3074 => 32759,
		3075 => 32759,
		3076 => 32759,
		3077 => 32759,
		3078 => 32759,
		3079 => 32759,
		3080 => 32759,
		3081 => 32759,
		3082 => 32759,
		3083 => 32759,
		3084 => 32759,
		3085 => 32759,
		3086 => 32759,
		3087 => 32759,
		3088 => 32759,
		3089 => 32759,
		3090 => 32759,
		3091 => 32759,
		3092 => 32759,
		3093 => 32759,
		3094 => 32759,
		3095 => 32759,
		3096 => 32759,
		3097 => 32759,
		3098 => 32759,
		3099 => 32759,
		3100 => 32759,
		3101 => 32759,
		3102 => 32759,
		3103 => 32759,
		3104 => 32759,
		3105 => 32759,
		3106 => 32759,
		3107 => 32759,
		3108 => 32759,
		3109 => 32759,
		3110 => 32759,
		3111 => 32759,
		3112 => 32759,
		3113 => 32759,
		3114 => 32759,
		3115 => 32759,
		3116 => 32759,
		3117 => 32759,
		3118 => 32759,
		3119 => 32759,
		3120 => 32759,
		3121 => 32760,
		3122 => 32760,
		3123 => 32760,
		3124 => 32760,
		3125 => 32760,
		3126 => 32760,
		3127 => 32760,
		3128 => 32760,
		3129 => 32760,
		3130 => 32760,
		3131 => 32760,
		3132 => 32760,
		3133 => 32760,
		3134 => 32760,
		3135 => 32760,
		3136 => 32760,
		3137 => 32760,
		3138 => 32760,
		3139 => 32760,
		3140 => 32760,
		3141 => 32760,
		3142 => 32760,
		3143 => 32760,
		3144 => 32760,
		3145 => 32760,
		3146 => 32760,
		3147 => 32760,
		3148 => 32760,
		3149 => 32760,
		3150 => 32760,
		3151 => 32760,
		3152 => 32760,
		3153 => 32760,
		3154 => 32760,
		3155 => 32760,
		3156 => 32760,
		3157 => 32760,
		3158 => 32760,
		3159 => 32760,
		3160 => 32760,
		3161 => 32760,
		3162 => 32760,
		3163 => 32760,
		3164 => 32760,
		3165 => 32760,
		3166 => 32760,
		3167 => 32760,
		3168 => 32760,
		3169 => 32760,
		3170 => 32760,
		3171 => 32760,
		3172 => 32760,
		3173 => 32760,
		3174 => 32761,
		3175 => 32761,
		3176 => 32761,
		3177 => 32761,
		3178 => 32761,
		3179 => 32761,
		3180 => 32761,
		3181 => 32761,
		3182 => 32761,
		3183 => 32761,
		3184 => 32761,
		3185 => 32761,
		3186 => 32761,
		3187 => 32761,
		3188 => 32761,
		3189 => 32761,
		3190 => 32761,
		3191 => 32761,
		3192 => 32761,
		3193 => 32761,
		3194 => 32761,
		3195 => 32761,
		3196 => 32761,
		3197 => 32761,
		3198 => 32761,
		3199 => 32761,
		3200 => 32761,
		3201 => 32761,
		3202 => 32761,
		3203 => 32761,
		3204 => 32761,
		3205 => 32761,
		3206 => 32761,
		3207 => 32761,
		3208 => 32761,
		3209 => 32761,
		3210 => 32761,
		3211 => 32761,
		3212 => 32761,
		3213 => 32761,
		3214 => 32761,
		3215 => 32761,
		3216 => 32761,
		3217 => 32761,
		3218 => 32761,
		3219 => 32761,
		3220 => 32761,
		3221 => 32761,
		3222 => 32761,
		3223 => 32761,
		3224 => 32761,
		3225 => 32761,
		3226 => 32761,
		3227 => 32761,
		3228 => 32761,
		3229 => 32761,
		3230 => 32761,
		3231 => 32761,
		3232 => 32761,
		3233 => 32761,
		3234 => 32761,
		3235 => 32761,
		3236 => 32762,
		3237 => 32762,
		3238 => 32762,
		3239 => 32762,
		3240 => 32762,
		3241 => 32762,
		3242 => 32762,
		3243 => 32762,
		3244 => 32762,
		3245 => 32762,
		3246 => 32762,
		3247 => 32762,
		3248 => 32762,
		3249 => 32762,
		3250 => 32762,
		3251 => 32762,
		3252 => 32762,
		3253 => 32762,
		3254 => 32762,
		3255 => 32762,
		3256 => 32762,
		3257 => 32762,
		3258 => 32762,
		3259 => 32762,
		3260 => 32762,
		3261 => 32762,
		3262 => 32762,
		3263 => 32762,
		3264 => 32762,
		3265 => 32762,
		3266 => 32762,
		3267 => 32762,
		3268 => 32762,
		3269 => 32762,
		3270 => 32762,
		3271 => 32762,
		3272 => 32762,
		3273 => 32762,
		3274 => 32762,
		3275 => 32762,
		3276 => 32762,
		3277 => 32762,
		3278 => 32762,
		3279 => 32762,
		3280 => 32762,
		3281 => 32762,
		3282 => 32762,
		3283 => 32762,
		3284 => 32762,
		3285 => 32762,
		3286 => 32762,
		3287 => 32762,
		3288 => 32762,
		3289 => 32762,
		3290 => 32762,
		3291 => 32762,
		3292 => 32762,
		3293 => 32762,
		3294 => 32762,
		3295 => 32762,
		3296 => 32762,
		3297 => 32762,
		3298 => 32762,
		3299 => 32762,
		3300 => 32762,
		3301 => 32762,
		3302 => 32762,
		3303 => 32762,
		3304 => 32762,
		3305 => 32762,
		3306 => 32762,
		3307 => 32762,
		3308 => 32762,
		3309 => 32762,
		3310 => 32762,
		3311 => 32763,
		3312 => 32763,
		3313 => 32763,
		3314 => 32763,
		3315 => 32763,
		3316 => 32763,
		3317 => 32763,
		3318 => 32763,
		3319 => 32763,
		3320 => 32763,
		3321 => 32763,
		3322 => 32763,
		3323 => 32763,
		3324 => 32763,
		3325 => 32763,
		3326 => 32763,
		3327 => 32763,
		3328 => 32763,
		3329 => 32763,
		3330 => 32763,
		3331 => 32763,
		3332 => 32763,
		3333 => 32763,
		3334 => 32763,
		3335 => 32763,
		3336 => 32763,
		3337 => 32763,
		3338 => 32763,
		3339 => 32763,
		3340 => 32763,
		3341 => 32763,
		3342 => 32763,
		3343 => 32763,
		3344 => 32763,
		3345 => 32763,
		3346 => 32763,
		3347 => 32763,
		3348 => 32763,
		3349 => 32763,
		3350 => 32763,
		3351 => 32763,
		3352 => 32763,
		3353 => 32763,
		3354 => 32763,
		3355 => 32763,
		3356 => 32763,
		3357 => 32763,
		3358 => 32763,
		3359 => 32763,
		3360 => 32763,
		3361 => 32763,
		3362 => 32763,
		3363 => 32763,
		3364 => 32763,
		3365 => 32763,
		3366 => 32763,
		3367 => 32763,
		3368 => 32763,
		3369 => 32763,
		3370 => 32763,
		3371 => 32763,
		3372 => 32763,
		3373 => 32763,
		3374 => 32763,
		3375 => 32763,
		3376 => 32763,
		3377 => 32763,
		3378 => 32763,
		3379 => 32763,
		3380 => 32763,
		3381 => 32763,
		3382 => 32763,
		3383 => 32763,
		3384 => 32763,
		3385 => 32763,
		3386 => 32763,
		3387 => 32763,
		3388 => 32763,
		3389 => 32763,
		3390 => 32763,
		3391 => 32763,
		3392 => 32763,
		3393 => 32763,
		3394 => 32763,
		3395 => 32763,
		3396 => 32763,
		3397 => 32763,
		3398 => 32763,
		3399 => 32763,
		3400 => 32763,
		3401 => 32763,
		3402 => 32763,
		3403 => 32763,
		3404 => 32763,
		3405 => 32764,
		3406 => 32764,
		3407 => 32764,
		3408 => 32764,
		3409 => 32764,
		3410 => 32764,
		3411 => 32764,
		3412 => 32764,
		3413 => 32764,
		3414 => 32764,
		3415 => 32764,
		3416 => 32764,
		3417 => 32764,
		3418 => 32764,
		3419 => 32764,
		3420 => 32764,
		3421 => 32764,
		3422 => 32764,
		3423 => 32764,
		3424 => 32764,
		3425 => 32764,
		3426 => 32764,
		3427 => 32764,
		3428 => 32764,
		3429 => 32764,
		3430 => 32764,
		3431 => 32764,
		3432 => 32764,
		3433 => 32764,
		3434 => 32764,
		3435 => 32764,
		3436 => 32764,
		3437 => 32764,
		3438 => 32764,
		3439 => 32764,
		3440 => 32764,
		3441 => 32764,
		3442 => 32764,
		3443 => 32764,
		3444 => 32764,
		3445 => 32764,
		3446 => 32764,
		3447 => 32764,
		3448 => 32764,
		3449 => 32764,
		3450 => 32764,
		3451 => 32764,
		3452 => 32764,
		3453 => 32764,
		3454 => 32764,
		3455 => 32764,
		3456 => 32764,
		3457 => 32764,
		3458 => 32764,
		3459 => 32764,
		3460 => 32764,
		3461 => 32764,
		3462 => 32764,
		3463 => 32764,
		3464 => 32764,
		3465 => 32764,
		3466 => 32764,
		3467 => 32764,
		3468 => 32764,
		3469 => 32764,
		3470 => 32764,
		3471 => 32764,
		3472 => 32764,
		3473 => 32764,
		3474 => 32764,
		3475 => 32764,
		3476 => 32764,
		3477 => 32764,
		3478 => 32764,
		3479 => 32764,
		3480 => 32764,
		3481 => 32764,
		3482 => 32764,
		3483 => 32764,
		3484 => 32764,
		3485 => 32764,
		3486 => 32764,
		3487 => 32764,
		3488 => 32764,
		3489 => 32764,
		3490 => 32764,
		3491 => 32764,
		3492 => 32764,
		3493 => 32764,
		3494 => 32764,
		3495 => 32764,
		3496 => 32764,
		3497 => 32764,
		3498 => 32764,
		3499 => 32764,
		3500 => 32764,
		3501 => 32764,
		3502 => 32764,
		3503 => 32764,
		3504 => 32764,
		3505 => 32764,
		3506 => 32764,
		3507 => 32764,
		3508 => 32764,
		3509 => 32764,
		3510 => 32764,
		3511 => 32764,
		3512 => 32764,
		3513 => 32764,
		3514 => 32764,
		3515 => 32764,
		3516 => 32764,
		3517 => 32764,
		3518 => 32764,
		3519 => 32764,
		3520 => 32764,
		3521 => 32764,
		3522 => 32764,
		3523 => 32764,
		3524 => 32764,
		3525 => 32764,
		3526 => 32764,
		3527 => 32764,
		3528 => 32764,
		3529 => 32764,
		3530 => 32765,
		3531 => 32765,
		3532 => 32765,
		3533 => 32765,
		3534 => 32765,
		3535 => 32765,
		3536 => 32765,
		3537 => 32765,
		3538 => 32765,
		3539 => 32765,
		3540 => 32765,
		3541 => 32765,
		3542 => 32765,
		3543 => 32765,
		3544 => 32765,
		3545 => 32765,
		3546 => 32765,
		3547 => 32765,
		3548 => 32765,
		3549 => 32765,
		3550 => 32765,
		3551 => 32765,
		3552 => 32765,
		3553 => 32765,
		3554 => 32765,
		3555 => 32765,
		3556 => 32765,
		3557 => 32765,
		3558 => 32765,
		3559 => 32765,
		3560 => 32765,
		3561 => 32765,
		3562 => 32765,
		3563 => 32765,
		3564 => 32765,
		3565 => 32765,
		3566 => 32765,
		3567 => 32765,
		3568 => 32765,
		3569 => 32765,
		3570 => 32765,
		3571 => 32765,
		3572 => 32765,
		3573 => 32765,
		3574 => 32765,
		3575 => 32765,
		3576 => 32765,
		3577 => 32765,
		3578 => 32765,
		3579 => 32765,
		3580 => 32765,
		3581 => 32765,
		3582 => 32765,
		3583 => 32765,
		3584 => 32765,
		3585 => 32765,
		3586 => 32765,
		3587 => 32765,
		3588 => 32765,
		3589 => 32765,
		3590 => 32765,
		3591 => 32765,
		3592 => 32765,
		3593 => 32765,
		3594 => 32765,
		3595 => 32765,
		3596 => 32765,
		3597 => 32765,
		3598 => 32765,
		3599 => 32765,
		3600 => 32765,
		3601 => 32765,
		3602 => 32765,
		3603 => 32765,
		3604 => 32765,
		3605 => 32765,
		3606 => 32765,
		3607 => 32765,
		3608 => 32765,
		3609 => 32765,
		3610 => 32765,
		3611 => 32765,
		3612 => 32765,
		3613 => 32765,
		3614 => 32765,
		3615 => 32765,
		3616 => 32765,
		3617 => 32765,
		3618 => 32765,
		3619 => 32765,
		3620 => 32765,
		3621 => 32765,
		3622 => 32765,
		3623 => 32765,
		3624 => 32765,
		3625 => 32765,
		3626 => 32765,
		3627 => 32765,
		3628 => 32765,
		3629 => 32765,
		3630 => 32765,
		3631 => 32765,
		3632 => 32765,
		3633 => 32765,
		3634 => 32765,
		3635 => 32765,
		3636 => 32765,
		3637 => 32765,
		3638 => 32765,
		3639 => 32765,
		3640 => 32765,
		3641 => 32765,
		3642 => 32765,
		3643 => 32765,
		3644 => 32765,
		3645 => 32765,
		3646 => 32765,
		3647 => 32765,
		3648 => 32765,
		3649 => 32765,
		3650 => 32765,
		3651 => 32765,
		3652 => 32765,
		3653 => 32765,
		3654 => 32765,
		3655 => 32765,
		3656 => 32765,
		3657 => 32765,
		3658 => 32765,
		3659 => 32765,
		3660 => 32765,
		3661 => 32765,
		3662 => 32765,
		3663 => 32765,
		3664 => 32765,
		3665 => 32765,
		3666 => 32765,
		3667 => 32765,
		3668 => 32765,
		3669 => 32765,
		3670 => 32765,
		3671 => 32765,
		3672 => 32765,
		3673 => 32765,
		3674 => 32765,
		3675 => 32765,
		3676 => 32765,
		3677 => 32765,
		3678 => 32765,
		3679 => 32765,
		3680 => 32765,
		3681 => 32765,
		3682 => 32765,
		3683 => 32765,
		3684 => 32765,
		3685 => 32765,
		3686 => 32765,
		3687 => 32765,
		3688 => 32765,
		3689 => 32765,
		3690 => 32765,
		3691 => 32765,
		3692 => 32765,
		3693 => 32765,
		3694 => 32765,
		3695 => 32765,
		3696 => 32765,
		3697 => 32765,
		3698 => 32765,
		3699 => 32765,
		3700 => 32765,
		3701 => 32765,
		3702 => 32765,
		3703 => 32765,
		3704 => 32765,
		3705 => 32765,
		3706 => 32765,
		3707 => 32765,
		3708 => 32765,
		3709 => 32765,
		3710 => 32765,
		3711 => 32765,
		3712 => 32765,
		3713 => 32765,
		3714 => 32765,
		3715 => 32765,
		3716 => 32765,
		3717 => 32765,
		3718 => 32765,
		3719 => 32765,
		3720 => 32766,
		3721 => 32766,
		3722 => 32766,
		3723 => 32766,
		3724 => 32766,
		3725 => 32766,
		3726 => 32766,
		3727 => 32766,
		3728 => 32766,
		3729 => 32766,
		3730 => 32766,
		3731 => 32766,
		3732 => 32766,
		3733 => 32766,
		3734 => 32766,
		3735 => 32766,
		3736 => 32766,
		3737 => 32766,
		3738 => 32766,
		3739 => 32766,
		3740 => 32766,
		3741 => 32766,
		3742 => 32766,
		3743 => 32766,
		3744 => 32766,
		3745 => 32766,
		3746 => 32766,
		3747 => 32766,
		3748 => 32766,
		3749 => 32766,
		3750 => 32766,
		3751 => 32766,
		3752 => 32766,
		3753 => 32766,
		3754 => 32766,
		3755 => 32766,
		3756 => 32766,
		3757 => 32766,
		3758 => 32766,
		3759 => 32766,
		3760 => 32766,
		3761 => 32766,
		3762 => 32766,
		3763 => 32766,
		3764 => 32766,
		3765 => 32766,
		3766 => 32766,
		3767 => 32766,
		3768 => 32766,
		3769 => 32766,
		3770 => 32766,
		3771 => 32766,
		3772 => 32766,
		3773 => 32766,
		3774 => 32766,
		3775 => 32766,
		3776 => 32766,
		3777 => 32766,
		3778 => 32766,
		3779 => 32766,
		3780 => 32766,
		3781 => 32766,
		3782 => 32766,
		3783 => 32766,
		3784 => 32766,
		3785 => 32766,
		3786 => 32766,
		3787 => 32766,
		3788 => 32766,
		3789 => 32766,
		3790 => 32766,
		3791 => 32766,
		3792 => 32766,
		3793 => 32766,
		3794 => 32766,
		3795 => 32766,
		3796 => 32766,
		3797 => 32766,
		3798 => 32766,
		3799 => 32766,
		3800 => 32766,
		3801 => 32766,
		3802 => 32766,
		3803 => 32766,
		3804 => 32766,
		3805 => 32766,
		3806 => 32766,
		3807 => 32766,
		3808 => 32766,
		3809 => 32766,
		3810 => 32766,
		3811 => 32766,
		3812 => 32766,
		3813 => 32766,
		3814 => 32766,
		3815 => 32766,
		3816 => 32766,
		3817 => 32766,
		3818 => 32766,
		3819 => 32766,
		3820 => 32766,
		3821 => 32766,
		3822 => 32766,
		3823 => 32766,
		3824 => 32766,
		3825 => 32766,
		3826 => 32766,
		3827 => 32766,
		3828 => 32766,
		3829 => 32766,
		3830 => 32766,
		3831 => 32766,
		3832 => 32766,
		3833 => 32766,
		3834 => 32766,
		3835 => 32766,
		3836 => 32766,
		3837 => 32766,
		3838 => 32766,
		3839 => 32766,
		3840 => 32766,
		3841 => 32766,
		3842 => 32766,
		3843 => 32766,
		3844 => 32766,
		3845 => 32766,
		3846 => 32766,
		3847 => 32766,
		3848 => 32766,
		3849 => 32766,
		3850 => 32766,
		3851 => 32766,
		3852 => 32766,
		3853 => 32766,
		3854 => 32766,
		3855 => 32766,
		3856 => 32766,
		3857 => 32766,
		3858 => 32766,
		3859 => 32766,
		3860 => 32766,
		3861 => 32766,
		3862 => 32766,
		3863 => 32766,
		3864 => 32766,
		3865 => 32766,
		3866 => 32766,
		3867 => 32766,
		3868 => 32766,
		3869 => 32766,
		3870 => 32766,
		3871 => 32766,
		3872 => 32766,
		3873 => 32766,
		3874 => 32766,
		3875 => 32766,
		3876 => 32766,
		3877 => 32766,
		3878 => 32766,
		3879 => 32766,
		3880 => 32766,
		3881 => 32766,
		3882 => 32766,
		3883 => 32766,
		3884 => 32766,
		3885 => 32766,
		3886 => 32766,
		3887 => 32766,
		3888 => 32766,
		3889 => 32766,
		3890 => 32766,
		3891 => 32766,
		3892 => 32766,
		3893 => 32766,
		3894 => 32766,
		3895 => 32766,
		3896 => 32766,
		3897 => 32766,
		3898 => 32766,
		3899 => 32766,
		3900 => 32766,
		3901 => 32766,
		3902 => 32766,
		3903 => 32766,
		3904 => 32766,
		3905 => 32766,
		3906 => 32766,
		3907 => 32766,
		3908 => 32766,
		3909 => 32766,
		3910 => 32766,
		3911 => 32766,
		3912 => 32766,
		3913 => 32766,
		3914 => 32766,
		3915 => 32766,
		3916 => 32766,
		3917 => 32766,
		3918 => 32766,
		3919 => 32766,
		3920 => 32766,
		3921 => 32766,
		3922 => 32766,
		3923 => 32766,
		3924 => 32766,
		3925 => 32766,
		3926 => 32766,
		3927 => 32766,
		3928 => 32766,
		3929 => 32766,
		3930 => 32766,
		3931 => 32766,
		3932 => 32766,
		3933 => 32766,
		3934 => 32766,
		3935 => 32766,
		3936 => 32766,
		3937 => 32766,
		3938 => 32766,
		3939 => 32766,
		3940 => 32766,
		3941 => 32766,
		3942 => 32766,
		3943 => 32766,
		3944 => 32766,
		3945 => 32766,
		3946 => 32766,
		3947 => 32766,
		3948 => 32766,
		3949 => 32766,
		3950 => 32766,
		3951 => 32766,
		3952 => 32766,
		3953 => 32766,
		3954 => 32766,
		3955 => 32766,
		3956 => 32766,
		3957 => 32766,
		3958 => 32766,
		3959 => 32766,
		3960 => 32766,
		3961 => 32766,
		3962 => 32766,
		3963 => 32766,
		3964 => 32766,
		3965 => 32766,
		3966 => 32766,
		3967 => 32766,
		3968 => 32766,
		3969 => 32766,
		3970 => 32766,
		3971 => 32766,
		3972 => 32766,
		3973 => 32766,
		3974 => 32766,
		3975 => 32766,
		3976 => 32766,
		3977 => 32766,
		3978 => 32766,
		3979 => 32766,
		3980 => 32766,
		3981 => 32766,
		3982 => 32766,
		3983 => 32766,
		3984 => 32766,
		3985 => 32766,
		3986 => 32766,
		3987 => 32766,
		3988 => 32766,
		3989 => 32766,
		3990 => 32766,
		3991 => 32766,
		3992 => 32766,
		3993 => 32766,
		3994 => 32766,
		3995 => 32766,
		3996 => 32766,
		3997 => 32766,
		3998 => 32766,
		3999 => 32766,
		4000 => 32766,
		4001 => 32766,
		4002 => 32766,
		4003 => 32766,
		4004 => 32766,
		4005 => 32766,
		4006 => 32766,
		4007 => 32766,
		4008 => 32766,
		4009 => 32766,
		4010 => 32766,
		4011 => 32766,
		4012 => 32766,
		4013 => 32766,
		4014 => 32766,
		4015 => 32766,
		4016 => 32766,
		4017 => 32766,
		4018 => 32766,
		4019 => 32766,
		4020 => 32766,
		4021 => 32766,
		4022 => 32766,
		4023 => 32766,
		4024 => 32766,
		4025 => 32766,
		4026 => 32766,
		4027 => 32766,
		4028 => 32766,
		4029 => 32766,
		4030 => 32766,
		4031 => 32766,
		4032 => 32766,
		4033 => 32766,
		4034 => 32766,
		4035 => 32766,
		4036 => 32766,
		4037 => 32766,
		4038 => 32766,
		4039 => 32766,
		4040 => 32766,
		4041 => 32766,
		4042 => 32766,
		4043 => 32766,
		4044 => 32766,
		4045 => 32766,
		4046 => 32766,
		4047 => 32766,
		4048 => 32766,
		4049 => 32766,
		4050 => 32766,
		4051 => 32766,
		4052 => 32766,
		4053 => 32766,
		4054 => 32766,
		4055 => 32766,
		4056 => 32766,
		4057 => 32766,
		4058 => 32766,
		4059 => 32766,
		4060 => 32766,
		4061 => 32766,
		4062 => 32766,
		4063 => 32766,
		4064 => 32766,
		4065 => 32766,
		4066 => 32766,
		4067 => 32766,
		4068 => 32766,
		4069 => 32766,
		4070 => 32766,
		4071 => 32766,
		4072 => 32766,
		4073 => 32766,
		4074 => 32766,
		4075 => 32766,
		4076 => 32766,
		4077 => 32766,
		4078 => 32766,
		4079 => 32766,
		4080 => 32766,
		4081 => 32766,
		4082 => 32766,
		4083 => 32766,
		4084 => 32766,
		4085 => 32766,
		4086 => 32766,
		4087 => 32766,
		4088 => 32766,
		4089 => 32766,
		4090 => 32766,
		4091 => 32766,
		4092 => 32766,
		4093 => 32766,
		4094 => 32766,
		4095 => 32766
);

begin
	dds_out <= std_logic_vector(TO_SIGNED(LUT(TO_INTEGER(unsigned(address))),16));
end beh;
